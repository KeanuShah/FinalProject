
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity Button_TenSec is
    port(clk, rst: in std_logic;
         addr: in std_logic_vector(9 downto 0);
         dout: out std_logic_vector(7 downto 0));
end Button_TenSec;

architecture Behavioral of Button_TenSec is

    type mem is array (0 to 951) of std_logic_vector(7 downto 0);
    signal Ten: mem := (
        0 => "00000001",
        1 => "00000001",
        2 => "00000001",
        3 => "00000001",
        4 => "00000000",
        5 => "00000000",
        6 => "00000000",
        7 => "00000000",
        8 => "00000000",
        9 => "00000000",
        10 => "00000000",
        11 => "00000000",
        12 => "00000000",
        13 => "00000000",
        14 => "00000000",
        15 => "00000000",
        16 => "00000000",
        17 => "00000000",
        18 => "00000000",
        19 => "00000000",
        20 => "00000000",
        21 => "00000000",
        22 => "00000000",
        23 => "00000000",
        24 => "00000000",
        25 => "00000000",
        26 => "00000000",
        27 => "00000000",
        28 => "00000000",
        29 => "00000000",
        30 => "00000000",
        31 => "00000001",
        32 => "00000001",
        33 => "00000001",
        34 => "00000001",
        35 => "00000001",
        36 => "00100101",
        37 => "10110111",
        38 => "11011111",
        39 => "11011111",
        40 => "11011111",
        41 => "11011111",
        42 => "11011111",
        43 => "11011111",
        44 => "11011111",
        45 => "11011111",
        46 => "11011111",
        47 => "11011111",
        48 => "11011111",
        49 => "11011111",
        50 => "11011111",
        51 => "11011111",
        52 => "11011111",
        53 => "11111111",
        54 => "11011111",
        55 => "11011111",
        56 => "11111111",
        57 => "11011111",
        58 => "11011111",
        59 => "11011111",
        60 => "11011111",
        61 => "11011111",
        62 => "11011111",
        63 => "11011111",
        64 => "10010111",
        65 => "00100101",
        66 => "00000001",
        67 => "00000001",
        68 => "00000001",
        69 => "00100001",
        70 => "11111111",
        71 => "11011111",
        72 => "11011111",
        73 => "11011111",
        74 => "11011111",
        75 => "11011111",
        76 => "11011111",
        77 => "11011111",
        78 => "11011111",
        79 => "11011110",
        80 => "11011110",
        81 => "11011111",
        82 => "11011111",
        83 => "11011111",
        84 => "11011111",
        85 => "11011111",
        86 => "11011111",
        87 => "11011111",
        88 => "11011111",
        89 => "11011111",
        90 => "11011111",
        91 => "11011111",
        92 => "11011111",
        93 => "11011111",
        94 => "11011111",
        95 => "11011111",
        96 => "11011111",
        97 => "11011111",
        98 => "11111111",
        99 => "11111111",
        100 => "00100101",
        101 => "00000001",
        102 => "00000000",
        103 => "10110011",
        104 => "11011111",
        105 => "10011010",
        106 => "00110000",
        107 => "00001100",
        108 => "00001100",
        109 => "00001100",
        110 => "00101100",
        111 => "00101100",
        112 => "00010000",
        113 => "00010000",
        114 => "00010000",
        115 => "00010000",
        116 => "00001100",
        117 => "00001100",
        118 => "00001100",
        119 => "00001100",
        120 => "00101100",
        121 => "00001100",
        122 => "00010000",
        123 => "00010000",
        124 => "00001100",
        125 => "00001100",
        126 => "00010000",
        127 => "00010000",
        128 => "00110000",
        129 => "00001100",
        130 => "00001100",
        131 => "00110000",
        132 => "10011010",
        133 => "11111111",
        134 => "10010011",
        135 => "00000001",
        136 => "00000000",
        137 => "11011111",
        138 => "11011111",
        139 => "00110000",
        140 => "00010000",
        141 => "00010000",
        142 => "00010000",
        143 => "00010000",
        144 => "00010000",
        145 => "00010000",
        146 => "00010000",
        147 => "00010000",
        148 => "00010000",
        149 => "00010000",
        150 => "00010000",
        151 => "00010000",
        152 => "00010000",
        153 => "00010000",
        154 => "00010000",
        155 => "00010000",
        156 => "00010000",
        157 => "00010000",
        158 => "00010000",
        159 => "00010000",
        160 => "00010000",
        161 => "00010000",
        162 => "00010000",
        163 => "00010000",
        164 => "00010000",
        165 => "00010000",
        166 => "00110000",
        167 => "11011111",
        168 => "11011111",
        169 => "00000001",
        170 => "00000000",
        171 => "11011111",
        172 => "11011111",
        173 => "00001100",
        174 => "00010000",
        175 => "00010000",
        176 => "00010000",
        177 => "00010000",
        178 => "00010000",
        179 => "00010000",
        180 => "00010000",
        181 => "00010000",
        182 => "00010000",
        183 => "00010000",
        184 => "00010000",
        185 => "00010000",
        186 => "00010000",
        187 => "00010000",
        188 => "00010000",
        189 => "00010000",
        190 => "00010000",
        191 => "00010000",
        192 => "00010000",
        193 => "00010000",
        194 => "00010000",
        195 => "00010000",
        196 => "00010000",
        197 => "00010000",
        198 => "00010000",
        199 => "00010000",
        200 => "00010000",
        201 => "11011111",
        202 => "11011111",
        203 => "00000000",
        204 => "00000000",
        205 => "11011111",
        206 => "11011111",
        207 => "00010000",
        208 => "00010000",
        209 => "00010000",
        210 => "00010000",
        211 => "00010000",
        212 => "00010000",
        213 => "00010000",
        214 => "00010000",
        215 => "00010000",
        216 => "00010000",
        217 => "00010000",
        218 => "00010000",
        219 => "00010000",
        220 => "00010000",
        221 => "00010000",
        222 => "00010000",
        223 => "00010000",
        224 => "00010000",
        225 => "00010000",
        226 => "00010000",
        227 => "00010000",
        228 => "00010000",
        229 => "00010000",
        230 => "00010000",
        231 => "00010000",
        232 => "00010000",
        233 => "00010000",
        234 => "00001100",
        235 => "11011111",
        236 => "11011111",
        237 => "00000000",
        238 => "00000000",
        239 => "11011111",
        240 => "11011111",
        241 => "00001100",
        242 => "00010000",
        243 => "00010000",
        244 => "00010000",
        245 => "00010000",
        246 => "00010000",
        247 => "00010000",
        248 => "00010000",
        249 => "00010000",
        250 => "00010000",
        251 => "00010000",
        252 => "00010000",
        253 => "00010000",
        254 => "00010000",
        255 => "00010000",
        256 => "00010000",
        257 => "00010000",
        258 => "00010000",
        259 => "00010000",
        260 => "00010000",
        261 => "00010000",
        262 => "00010000",
        263 => "00010000",
        264 => "00010000",
        265 => "00010000",
        266 => "00010000",
        267 => "00010000",
        268 => "00010000",
        269 => "11011111",
        270 => "11011111",
        271 => "00000000",
        272 => "00000000",
        273 => "11111111",
        274 => "11011111",
        275 => "00010000",
        276 => "00010000",
        277 => "00010000",
        278 => "00010000",
        279 => "00010000",
        280 => "00010000",
        281 => "00010000",
        282 => "00010000",
        283 => "00010000",
        284 => "00010000",
        285 => "00010000",
        286 => "00010000",
        287 => "00010000",
        288 => "00010000",
        289 => "00010000",
        290 => "00010000",
        291 => "00010100",
        292 => "00010000",
        293 => "00010000",
        294 => "00010100",
        295 => "00010000",
        296 => "00010000",
        297 => "00010000",
        298 => "00010000",
        299 => "00010000",
        300 => "00010000",
        301 => "00010000",
        302 => "00010000",
        303 => "10111111",
        304 => "11011111",
        305 => "00000000",
        306 => "00000000",
        307 => "11111111",
        308 => "11011111",
        309 => "00010000",
        310 => "00010000",
        311 => "00010000",
        312 => "00010000",
        313 => "00010000",
        314 => "00010000",
        315 => "00010000",
        316 => "00010000",
        317 => "00010000",
        318 => "00010000",
        319 => "00010000",
        320 => "00010000",
        321 => "00010000",
        322 => "00010000",
        323 => "00010000",
        324 => "00010000",
        325 => "00010000",
        326 => "00010000",
        327 => "00010100",
        328 => "00010000",
        329 => "00010100",
        330 => "00010000",
        331 => "00010100",
        332 => "00010000",
        333 => "00010100",
        334 => "00010000",
        335 => "00010000",
        336 => "00010000",
        337 => "10111111",
        338 => "11011111",
        339 => "00000000",
        340 => "00000000",
        341 => "11111111",
        342 => "11011111",
        343 => "00101100",
        344 => "00010000",
        345 => "00010000",
        346 => "00010000",
        347 => "00010000",
        348 => "00010000",
        349 => "00110101",
        350 => "10111110",
        351 => "10111110",
        352 => "00010000",
        353 => "00010000",
        354 => "00010000",
        355 => "01111101",
        356 => "10111110",
        357 => "11011110",
        358 => "11011110",
        359 => "01010100",
        360 => "00010000",
        361 => "00010000",
        362 => "00010000",
        363 => "00010000",
        364 => "00010000",
        365 => "00010000",
        366 => "00010000",
        367 => "00010000",
        368 => "00010100",
        369 => "00010000",
        370 => "00001100",
        371 => "11011111",
        372 => "11011111",
        373 => "00000000",
        374 => "00000000",
        375 => "11111111",
        376 => "11011111",
        377 => "00101100",
        378 => "00010000",
        379 => "00010000",
        380 => "00010000",
        381 => "00010000",
        382 => "00111001",
        383 => "10111111",
        384 => "11011110",
        385 => "11011110",
        386 => "00010000",
        387 => "00010000",
        388 => "00110101",
        389 => "10111111",
        390 => "01110101",
        391 => "01001100",
        392 => "11011010",
        393 => "11011110",
        394 => "00010000",
        395 => "00010000",
        396 => "00010000",
        397 => "00010000",
        398 => "00010000",
        399 => "00010000",
        400 => "00010000",
        401 => "00010000",
        402 => "00010000",
        403 => "00010000",
        404 => "00010000",
        405 => "11011111",
        406 => "11011111",
        407 => "00000000",
        408 => "00000000",
        409 => "11011111",
        410 => "11011111",
        411 => "00010000",
        412 => "00010000",
        413 => "00010000",
        414 => "00010000",
        415 => "00010000",
        416 => "10011110",
        417 => "01111010",
        418 => "10111110",
        419 => "10111110",
        420 => "00010000",
        421 => "00010000",
        422 => "10011110",
        423 => "10111110",
        424 => "01010001",
        425 => "00110001",
        426 => "11011111",
        427 => "11011111",
        428 => "01010100",
        429 => "00110000",
        430 => "10111101",
        431 => "11011110",
        432 => "10111110",
        433 => "10111110",
        434 => "00010100",
        435 => "00010000",
        436 => "00010100",
        437 => "00010000",
        438 => "00101100",
        439 => "11011111",
        440 => "11111111",
        441 => "00000000",
        442 => "00000000",
        443 => "11011111",
        444 => "11011111",
        445 => "00010000",
        446 => "00010000",
        447 => "00010000",
        448 => "00010000",
        449 => "00010000",
        450 => "00010000",
        451 => "00110000",
        452 => "10111110",
        453 => "10111110",
        454 => "00010000",
        455 => "00010000",
        456 => "10111110",
        457 => "10111110",
        458 => "00110000",
        459 => "10111110",
        460 => "10111010",
        461 => "11011111",
        462 => "01110101",
        463 => "10011001",
        464 => "11011110",
        465 => "01110001",
        466 => "00101100",
        467 => "00101100",
        468 => "00010000",
        469 => "00010000",
        470 => "00010000",
        471 => "00010000",
        472 => "00001100",
        473 => "11011111",
        474 => "11111111",
        475 => "00000000",
        476 => "00000000",
        477 => "11011111",
        478 => "11011111",
        479 => "00010000",
        480 => "00010000",
        481 => "00010000",
        482 => "00010000",
        483 => "00010000",
        484 => "00010000",
        485 => "00010000",
        486 => "10111110",
        487 => "10111110",
        488 => "00010000",
        489 => "00010000",
        490 => "10111110",
        491 => "11011110",
        492 => "10111110",
        493 => "10011001",
        494 => "01110101",
        495 => "10111111",
        496 => "01111001",
        497 => "01110100",
        498 => "11011110",
        499 => "11011111",
        500 => "10111110",
        501 => "00101100",
        502 => "00010000",
        503 => "00010000",
        504 => "00010000",
        505 => "00010000",
        506 => "00010000",
        507 => "11011111",
        508 => "11011111",
        509 => "00000000",
        510 => "00000000",
        511 => "11011111",
        512 => "11011111",
        513 => "00010000",
        514 => "00010000",
        515 => "00010000",
        516 => "00010000",
        517 => "00010000",
        518 => "00010000",
        519 => "00010000",
        520 => "10111110",
        521 => "11011110",
        522 => "00010000",
        523 => "00010000",
        524 => "10011110",
        525 => "11011111",
        526 => "10011001",
        527 => "00101100",
        528 => "10011001",
        529 => "10111110",
        530 => "01010100",
        531 => "00001100",
        532 => "00101100",
        533 => "10111110",
        534 => "11011110",
        535 => "11011110",
        536 => "01111000",
        537 => "00010000",
        538 => "00010000",
        539 => "00010000",
        540 => "00010000",
        541 => "11011111",
        542 => "11011111",
        543 => "00000000",
        544 => "00000000",
        545 => "11011111",
        546 => "11011111",
        547 => "00001100",
        548 => "00010000",
        549 => "00010000",
        550 => "00010000",
        551 => "00010000",
        552 => "00010000",
        553 => "00101100",
        554 => "10111110",
        555 => "11011110",
        556 => "00101100",
        557 => "00001100",
        558 => "01010101",
        559 => "10111111",
        560 => "10011001",
        561 => "01001100",
        562 => "11011110",
        563 => "10111110",
        564 => "00010000",
        565 => "00010000",
        566 => "00001100",
        567 => "00101100",
        568 => "01110101",
        569 => "10111110",
        570 => "01111101",
        571 => "00010000",
        572 => "00010000",
        573 => "00010000",
        574 => "00010000",
        575 => "10111111",
        576 => "11011111",
        577 => "00000000",
        578 => "00000000",
        579 => "11011111",
        580 => "11011111",
        581 => "00001100",
        582 => "00010000",
        583 => "00010000",
        584 => "00010000",
        585 => "00010000",
        586 => "01111101",
        587 => "10111110",
        588 => "11011110",
        589 => "11011110",
        590 => "11011110",
        591 => "01111001",
        592 => "00010000",
        593 => "01111101",
        594 => "10111110",
        595 => "11011110",
        596 => "11011110",
        597 => "01010000",
        598 => "00010000",
        599 => "01111101",
        600 => "10111110",
        601 => "10111110",
        602 => "10111110",
        603 => "10011110",
        604 => "00010000",
        605 => "00010000",
        606 => "00010000",
        607 => "00010000",
        608 => "00001100",
        609 => "10111111",
        610 => "11011111",
        611 => "00000000",
        612 => "00000000",
        613 => "11011111",
        614 => "11011111",
        615 => "00010000",
        616 => "00010000",
        617 => "00010000",
        618 => "00010000",
        619 => "00010000",
        620 => "00010000",
        621 => "00010000",
        622 => "00010000",
        623 => "00010000",
        624 => "00010000",
        625 => "00010000",
        626 => "00010000",
        627 => "00010000",
        628 => "00010000",
        629 => "00010000",
        630 => "00010000",
        631 => "00010000",
        632 => "00010000",
        633 => "00010000",
        634 => "00010000",
        635 => "00010000",
        636 => "00010000",
        637 => "00010000",
        638 => "00010000",
        639 => "00010000",
        640 => "00010000",
        641 => "00010000",
        642 => "00010000",
        643 => "11011111",
        644 => "11011111",
        645 => "00000000",
        646 => "00000000",
        647 => "11011111",
        648 => "11011111",
        649 => "00001100",
        650 => "00010000",
        651 => "00010000",
        652 => "00010000",
        653 => "00010100",
        654 => "00010000",
        655 => "00010100",
        656 => "00010000",
        657 => "00010000",
        658 => "00010000",
        659 => "00010000",
        660 => "00010000",
        661 => "00010000",
        662 => "00010000",
        663 => "00010000",
        664 => "00010000",
        665 => "00010000",
        666 => "00010000",
        667 => "00010000",
        668 => "00010000",
        669 => "00010000",
        670 => "00010000",
        671 => "00010000",
        672 => "00010000",
        673 => "00010000",
        674 => "00010000",
        675 => "00010000",
        676 => "00010000",
        677 => "11011110",
        678 => "11011111",
        679 => "00000000",
        680 => "00000000",
        681 => "11011111",
        682 => "11011111",
        683 => "00010000",
        684 => "00010000",
        685 => "00010000",
        686 => "00010000",
        687 => "00010100",
        688 => "00010100",
        689 => "00010000",
        690 => "00010000",
        691 => "00010000",
        692 => "00010000",
        693 => "00010000",
        694 => "00010000",
        695 => "00010000",
        696 => "00010000",
        697 => "00010000",
        698 => "00010000",
        699 => "00010000",
        700 => "00010000",
        701 => "00010000",
        702 => "00010000",
        703 => "00010000",
        704 => "00010000",
        705 => "00010100",
        706 => "00010000",
        707 => "00010000",
        708 => "00010000",
        709 => "00010000",
        710 => "00010000",
        711 => "11011110",
        712 => "11011111",
        713 => "00000000",
        714 => "00000000",
        715 => "11111111",
        716 => "11011111",
        717 => "00010000",
        718 => "00010000",
        719 => "00010000",
        720 => "00010000",
        721 => "00010000",
        722 => "00010000",
        723 => "00010000",
        724 => "00010100",
        725 => "00010000",
        726 => "00010000",
        727 => "00010000",
        728 => "00010000",
        729 => "00010000",
        730 => "00010000",
        731 => "00010000",
        732 => "00010000",
        733 => "00010000",
        734 => "00010000",
        735 => "00010000",
        736 => "00010000",
        737 => "00010000",
        738 => "00010000",
        739 => "00010000",
        740 => "00010000",
        741 => "00010000",
        742 => "00010000",
        743 => "00010000",
        744 => "00010000",
        745 => "11011111",
        746 => "11011111",
        747 => "00000000",
        748 => "00000000",
        749 => "11111111",
        750 => "11011111",
        751 => "00010000",
        752 => "00010000",
        753 => "00010000",
        754 => "00010000",
        755 => "00010000",
        756 => "00010000",
        757 => "00010000",
        758 => "00010000",
        759 => "00010000",
        760 => "00010100",
        761 => "00010100",
        762 => "00010000",
        763 => "00010000",
        764 => "00010100",
        765 => "00010000",
        766 => "00010000",
        767 => "00010000",
        768 => "00010000",
        769 => "00010000",
        770 => "00010100",
        771 => "00010000",
        772 => "00010100",
        773 => "00010000",
        774 => "00010000",
        775 => "00010000",
        776 => "00010000",
        777 => "00010000",
        778 => "00001100",
        779 => "11011111",
        780 => "11011111",
        781 => "00000000",
        782 => "00000000",
        783 => "11111111",
        784 => "11011111",
        785 => "00101100",
        786 => "00010000",
        787 => "00010000",
        788 => "00010000",
        789 => "00010000",
        790 => "00010000",
        791 => "00010000",
        792 => "00010000",
        793 => "00010000",
        794 => "00010000",
        795 => "00010000",
        796 => "00010000",
        797 => "00010000",
        798 => "00010000",
        799 => "00010000",
        800 => "00010000",
        801 => "00010000",
        802 => "00010000",
        803 => "00010000",
        804 => "00010000",
        805 => "00010000",
        806 => "00010000",
        807 => "00010000",
        808 => "00010000",
        809 => "00010000",
        810 => "00010000",
        811 => "00010000",
        812 => "00110000",
        813 => "11011111",
        814 => "11011111",
        815 => "00000000",
        816 => "00000000",
        817 => "10110111",
        818 => "11011111",
        819 => "10011010",
        820 => "00101100",
        821 => "00101100",
        822 => "00101100",
        823 => "00001100",
        824 => "00001100",
        825 => "00001100",
        826 => "00001100",
        827 => "00010000",
        828 => "00010000",
        829 => "00010000",
        830 => "00010000",
        831 => "00001100",
        832 => "00010000",
        833 => "00001100",
        834 => "00001100",
        835 => "00001100",
        836 => "00010000",
        837 => "00010000",
        838 => "00001100",
        839 => "00001100",
        840 => "00001100",
        841 => "00001100",
        842 => "00001100",
        843 => "00110000",
        844 => "00001100",
        845 => "00110000",
        846 => "10011010",
        847 => "11011111",
        848 => "10010011",
        849 => "00000001",
        850 => "00000001",
        851 => "00000001",
        852 => "11011111",
        853 => "11011111",
        854 => "11011111",
        855 => "11011111",
        856 => "11011111",
        857 => "11011111",
        858 => "11011111",
        859 => "11011111",
        860 => "11011111",
        861 => "11011111",
        862 => "11011111",
        863 => "11011111",
        864 => "11011111",
        865 => "11011111",
        866 => "11011111",
        867 => "11011111",
        868 => "11011111",
        869 => "11011111",
        870 => "11011111",
        871 => "11011111",
        872 => "11011111",
        873 => "11011111",
        874 => "11011111",
        875 => "11011111",
        876 => "11011110",
        877 => "11011111",
        878 => "11011111",
        879 => "11011111",
        880 => "11111111",
        881 => "11011111",
        882 => "00100101",
        883 => "00000001",
        884 => "00000001",
        885 => "00000001",
        886 => "00000101",
        887 => "10010111",
        888 => "11011011",
        889 => "11011111",
        890 => "11111111",
        891 => "11011111",
        892 => "11011111",
        893 => "11011111",
        894 => "11011111",
        895 => "11011111",
        896 => "11111111",
        897 => "11111111",
        898 => "11111111",
        899 => "11111111",
        900 => "11111111",
        901 => "11011111",
        902 => "11111111",
        903 => "11011111",
        904 => "11011111",
        905 => "11011111",
        906 => "11011111",
        907 => "11011111",
        908 => "11011111",
        909 => "11011111",
        910 => "11011111",
        911 => "11011111",
        912 => "11011111",
        913 => "11011111",
        914 => "10010011",
        915 => "00100101",
        916 => "00000001",
        917 => "00000001",
        918 => "00000001",
        919 => "00000001",
        920 => "00000001",
        921 => "00000001",
        922 => "00000000",
        923 => "00000000",
        924 => "00000000",
        925 => "00000000",
        926 => "00000000",
        927 => "00000000",
        928 => "00000000",
        929 => "00000000",
        930 => "00000000",
        931 => "00000000",
        932 => "00000000",
        933 => "00000000",
        934 => "00000000",
        935 => "00000000",
        936 => "00000000",
        937 => "00000000",
        938 => "00000000",
        939 => "00000000",
        940 => "00000000",
        941 => "00000000",
        942 => "00000000",
        943 => "00000000",
        944 => "00000000",
        945 => "00000000",
        946 => "00000000",
        947 => "00000000",
        948 => "00000001",
        949 => "00000001",
        950 => "00000001",
        951 => "00000001");
begin

    process(clk)
    begin
    
        if rising_edge(clk) then
            if rst = '1' then
                Ten <= (others => (others => '0'));
            else
                dout <= Ten(to_integer(unsigned(addr)));
            end if;
        end if;
    end process;

end Behavioral;


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity Button_TwoSec is
    port(clk, rst: in std_logic;
             addr: in std_logic_vector(9 downto 0);
             dout: out std_logic_vector(7 downto 0));
end Button_TwoSec;

architecture Behavioral of Button_TwoSec is

     type mem is array (0 to 755) of std_logic_vector(7 downto 0);
     signal Two: mem := (
        0 => "00000001",
        1 => "00000001",
        2 => "00000001",
        3 => "00000001",
        4 => "00000000",
        5 => "00000000",
        6 => "00000000",
        7 => "00000000",
        8 => "00000000",
        9 => "00000000",
        10 => "00000000",
        11 => "00000000",
        12 => "00000000",
        13 => "00000000",
        14 => "00000000",
        15 => "00000000",
        16 => "00000000",
        17 => "00000000",
        18 => "00000000",
        19 => "00000000",
        20 => "00000000",
        21 => "00000000",
        22 => "00000000",
        23 => "00000000",
        24 => "00000001",
        25 => "00000001",
        26 => "00000001",
        27 => "00000001",
        28 => "00000001",
        29 => "00100101",
        30 => "10010111",
        31 => "11011111",
        32 => "11011111",
        33 => "11011111",
        34 => "11011111",
        35 => "11011111",
        36 => "11011111",
        37 => "11111111",
        38 => "11111111",
        39 => "11011111",
        40 => "11011111",
        41 => "11011111",
        42 => "11111111",
        43 => "11111111",
        44 => "11011111",
        45 => "11011111",
        46 => "11011111",
        47 => "11011111",
        48 => "11011111",
        49 => "11011011",
        50 => "10110111",
        51 => "00100101",
        52 => "00000001",
        53 => "00000001",
        54 => "00000001",
        55 => "00100101",
        56 => "11111111",
        57 => "11011111",
        58 => "11011111",
        59 => "11011111",
        60 => "11011111",
        61 => "11011111",
        62 => "11011111",
        63 => "11011111",
        64 => "11011111",
        65 => "11011111",
        66 => "11011111",
        67 => "11011111",
        68 => "11011111",
        69 => "11011111",
        70 => "11011111",
        71 => "11011111",
        72 => "11011111",
        73 => "11011111",
        74 => "11011111",
        75 => "11011111",
        76 => "11011111",
        77 => "11011111",
        78 => "11011111",
        79 => "00100101",
        80 => "00000001",
        81 => "00000001",
        82 => "10010011",
        83 => "11011111",
        84 => "10011010",
        85 => "00110000",
        86 => "00001100",
        87 => "00001100",
        88 => "00001100",
        89 => "00101100",
        90 => "00001100",
        91 => "00001100",
        92 => "00010000",
        93 => "00010000",
        94 => "00010000",
        95 => "00010000",
        96 => "00010000",
        97 => "00001100",
        98 => "00010000",
        99 => "00001100",
        100 => "00001100",
        101 => "00010000",
        102 => "00001100",
        103 => "00110000",
        104 => "10011010",
        105 => "11011111",
        106 => "10010011",
        107 => "00000001",
        108 => "00000000",
        109 => "11011111",
        110 => "11011111",
        111 => "00110000",
        112 => "00010000",
        113 => "00010000",
        114 => "00010000",
        115 => "00010000",
        116 => "00010000",
        117 => "00010000",
        118 => "00010000",
        119 => "00010000",
        120 => "00010000",
        121 => "00010000",
        122 => "00010000",
        123 => "00010000",
        124 => "00010000",
        125 => "00010000",
        126 => "00010000",
        127 => "00010000",
        128 => "00010000",
        129 => "00010000",
        130 => "00010000",
        131 => "00110000",
        132 => "11011111",
        133 => "11111111",
        134 => "00000000",
        135 => "00000000",
        136 => "11111111",
        137 => "11011111",
        138 => "00001100",
        139 => "00010000",
        140 => "00010000",
        141 => "00010000",
        142 => "00010000",
        143 => "00010000",
        144 => "00010000",
        145 => "00010000",
        146 => "00010000",
        147 => "00010000",
        148 => "00010000",
        149 => "00010000",
        150 => "00010000",
        151 => "00010000",
        152 => "00010000",
        153 => "00010000",
        154 => "00010000",
        155 => "00010000",
        156 => "00010100",
        157 => "00010000",
        158 => "00010000",
        159 => "11011111",
        160 => "11011111",
        161 => "00000000",
        162 => "00000000",
        163 => "11011111",
        164 => "11011111",
        165 => "00010000",
        166 => "00010000",
        167 => "00010000",
        168 => "00010100",
        169 => "00010000",
        170 => "00010000",
        171 => "00010000",
        172 => "00010000",
        173 => "00010000",
        174 => "00010000",
        175 => "00010000",
        176 => "00010000",
        177 => "00010000",
        178 => "00010000",
        179 => "00010000",
        180 => "00010000",
        181 => "00010000",
        182 => "00010000",
        183 => "00010000",
        184 => "00010000",
        185 => "00010000",
        186 => "11011111",
        187 => "11111111",
        188 => "00000001",
        189 => "00000000",
        190 => "11111111",
        191 => "11011111",
        192 => "00010000",
        193 => "00010000",
        194 => "00010000",
        195 => "00010000",
        196 => "00010000",
        197 => "00010000",
        198 => "00010000",
        199 => "00010000",
        200 => "00010000",
        201 => "00010000",
        202 => "00010000",
        203 => "00010000",
        204 => "00010000",
        205 => "00010000",
        206 => "00010000",
        207 => "00010000",
        208 => "00010000",
        209 => "00010000",
        210 => "00010000",
        211 => "00010000",
        212 => "00010000",
        213 => "11011111",
        214 => "11111111",
        215 => "00000001",
        216 => "00000000",
        217 => "11011111",
        218 => "11011111",
        219 => "00010000",
        220 => "00010000",
        221 => "00010000",
        222 => "00010000",
        223 => "00010000",
        224 => "00010000",
        225 => "00010000",
        226 => "00010100",
        227 => "00010100",
        228 => "00010000",
        229 => "00010000",
        230 => "00010000",
        231 => "00010000",
        232 => "00010000",
        233 => "00010000",
        234 => "00010000",
        235 => "00010000",
        236 => "00010000",
        237 => "00010000",
        238 => "00010000",
        239 => "00010000",
        240 => "11011111",
        241 => "11111111",
        242 => "00000001",
        243 => "00000000",
        244 => "11111111",
        245 => "11011111",
        246 => "00001100",
        247 => "00010000",
        248 => "00010000",
        249 => "00010000",
        250 => "00010000",
        251 => "00010000",
        252 => "00010000",
        253 => "00010000",
        254 => "00010000",
        255 => "00010000",
        256 => "00010000",
        257 => "00010000",
        258 => "00010000",
        259 => "00010000",
        260 => "00010000",
        261 => "00010000",
        262 => "00010000",
        263 => "00010000",
        264 => "00010000",
        265 => "00010100",
        266 => "00010000",
        267 => "11011111",
        268 => "11111111",
        269 => "00000001",
        270 => "00000000",
        271 => "11011111",
        272 => "11011111",
        273 => "00010000",
        274 => "00010000",
        275 => "00010000",
        276 => "00010000",
        277 => "00010000",
        278 => "10111110",
        279 => "11011110",
        280 => "10111110",
        281 => "10011110",
        282 => "00010000",
        283 => "00010000",
        284 => "00010000",
        285 => "00010000",
        286 => "00010000",
        287 => "00010000",
        288 => "00010000",
        289 => "00010100",
        290 => "00010000",
        291 => "00010100",
        292 => "00010000",
        293 => "00010000",
        294 => "11011111",
        295 => "11111111",
        296 => "00000001",
        297 => "00000000",
        298 => "11111111",
        299 => "11011111",
        300 => "00010000",
        301 => "00010000",
        302 => "00010000",
        303 => "00010100",
        304 => "00111000",
        305 => "10111110",
        306 => "01010000",
        307 => "01010001",
        308 => "10111111",
        309 => "01111001",
        310 => "00010000",
        311 => "00010000",
        312 => "00010000",
        313 => "00010000",
        314 => "00010000",
        315 => "00010000",
        316 => "00010000",
        317 => "00010000",
        318 => "00010000",
        319 => "00010000",
        320 => "00010000",
        321 => "11011111",
        322 => "11111111",
        323 => "00000001",
        324 => "00000000",
        325 => "11111111",
        326 => "11011111",
        327 => "00010000",
        328 => "00010000",
        329 => "00010000",
        330 => "00010000",
        331 => "00010000",
        332 => "00010000",
        333 => "00010000",
        334 => "00110001",
        335 => "10111111",
        336 => "10111101",
        337 => "00101100",
        338 => "00110000",
        339 => "10011110",
        340 => "10111110",
        341 => "10111110",
        342 => "10111101",
        343 => "00110100",
        344 => "00010000",
        345 => "00010000",
        346 => "00010000",
        347 => "00010000",
        348 => "11011111",
        349 => "11111111",
        350 => "00000001",
        351 => "00000000",
        352 => "11111111",
        353 => "11011111",
        354 => "00001100",
        355 => "00010000",
        356 => "00010000",
        357 => "00010000",
        358 => "00010000",
        359 => "00010000",
        360 => "00010000",
        361 => "00110101",
        362 => "10111111",
        363 => "01111001",
        364 => "00110000",
        365 => "01111001",
        366 => "10111110",
        367 => "01010001",
        368 => "00101100",
        369 => "00101100",
        370 => "00010000",
        371 => "00010000",
        372 => "00010000",
        373 => "00010000",
        374 => "00010000",
        375 => "11011111",
        376 => "11111111",
        377 => "00000001",
        378 => "00000000",
        379 => "11011111",
        380 => "11011111",
        381 => "00010000",
        382 => "00010000",
        383 => "00010000",
        384 => "00010000",
        385 => "00010000",
        386 => "00010000",
        387 => "00010000",
        388 => "10111110",
        389 => "10111110",
        390 => "00010000",
        391 => "00010000",
        392 => "00110101",
        393 => "10111111",
        394 => "11011111",
        395 => "11011110",
        396 => "00101100",
        397 => "00010000",
        398 => "00010000",
        399 => "00010000",
        400 => "00010000",
        401 => "00010000",
        402 => "11011111",
        403 => "11111111",
        404 => "00000001",
        405 => "00000000",
        406 => "11011111",
        407 => "11011111",
        408 => "00010000",
        409 => "00010000",
        410 => "00010000",
        411 => "00010000",
        412 => "00010000",
        413 => "00010000",
        414 => "10111110",
        415 => "10111110",
        416 => "00101100",
        417 => "00010000",
        418 => "00010000",
        419 => "00010000",
        420 => "00001100",
        421 => "10111110",
        422 => "11011110",
        423 => "11011110",
        424 => "01111000",
        425 => "00010000",
        426 => "00010000",
        427 => "00010000",
        428 => "00010000",
        429 => "11011111",
        430 => "11111111",
        431 => "00000001",
        432 => "00000000",
        433 => "11011111",
        434 => "11011111",
        435 => "00010000",
        436 => "00010000",
        437 => "00010000",
        438 => "00010000",
        439 => "00010000",
        440 => "10111110",
        441 => "10111110",
        442 => "01010000",
        443 => "00101100",
        444 => "00110000",
        445 => "00010000",
        446 => "00010000",
        447 => "00001100",
        448 => "00101100",
        449 => "01010101",
        450 => "11011110",
        451 => "10011101",
        452 => "00010000",
        453 => "00010000",
        454 => "00010000",
        455 => "00010000",
        456 => "11011111",
        457 => "11111111",
        458 => "00000001",
        459 => "00000000",
        460 => "11111111",
        461 => "10111111",
        462 => "00010000",
        463 => "00010100",
        464 => "00010000",
        465 => "00010000",
        466 => "01111101",
        467 => "10111110",
        468 => "11011110",
        469 => "11011110",
        470 => "10111110",
        471 => "10111101",
        472 => "00110100",
        473 => "01111101",
        474 => "10111110",
        475 => "10111110",
        476 => "10111110",
        477 => "10111101",
        478 => "00001100",
        479 => "00010000",
        480 => "00010000",
        481 => "00010000",
        482 => "00010000",
        483 => "11011111",
        484 => "11111111",
        485 => "00000001",
        486 => "00000000",
        487 => "11011111",
        488 => "10111111",
        489 => "00010000",
        490 => "00010000",
        491 => "00010000",
        492 => "00010000",
        493 => "00010000",
        494 => "00010000",
        495 => "00010000",
        496 => "00010000",
        497 => "00010000",
        498 => "00010000",
        499 => "00010000",
        500 => "00010000",
        501 => "00010000",
        502 => "00010000",
        503 => "00010000",
        504 => "00010000",
        505 => "00010000",
        506 => "00010000",
        507 => "00010100",
        508 => "00010000",
        509 => "00010000",
        510 => "11011111",
        511 => "11111111",
        512 => "00000001",
        513 => "00000000",
        514 => "11011111",
        515 => "11011111",
        516 => "00010000",
        517 => "00010000",
        518 => "00010000",
        519 => "00010000",
        520 => "00010000",
        521 => "00010000",
        522 => "00010000",
        523 => "00010000",
        524 => "00010000",
        525 => "00010000",
        526 => "00010000",
        527 => "00010000",
        528 => "00010000",
        529 => "00010000",
        530 => "00010000",
        531 => "00010000",
        532 => "00010000",
        533 => "00010000",
        534 => "00010100",
        535 => "00010000",
        536 => "00010000",
        537 => "11011111",
        538 => "11111111",
        539 => "00000001",
        540 => "00000000",
        541 => "11011111",
        542 => "11011111",
        543 => "00010000",
        544 => "00010000",
        545 => "00010000",
        546 => "00010000",
        547 => "00010000",
        548 => "00010000",
        549 => "00010000",
        550 => "00010000",
        551 => "00010000",
        552 => "00010000",
        553 => "00010000",
        554 => "00010000",
        555 => "00010000",
        556 => "00010000",
        557 => "00010100",
        558 => "00010000",
        559 => "00010000",
        560 => "00010000",
        561 => "00010100",
        562 => "00010000",
        563 => "00010000",
        564 => "11011111",
        565 => "11111111",
        566 => "00000001",
        567 => "00000000",
        568 => "11111111",
        569 => "11011111",
        570 => "00001100",
        571 => "00010000",
        572 => "00010000",
        573 => "00010100",
        574 => "00010000",
        575 => "00010000",
        576 => "00010000",
        577 => "00010000",
        578 => "00010100",
        579 => "00010000",
        580 => "00010000",
        581 => "00010000",
        582 => "00010000",
        583 => "00010000",
        584 => "00010000",
        585 => "00010000",
        586 => "00010000",
        587 => "00010000",
        588 => "00010000",
        589 => "00010000",
        590 => "00010000",
        591 => "11011111",
        592 => "11111111",
        593 => "00000001",
        594 => "00000000",
        595 => "11111111",
        596 => "11011111",
        597 => "00010000",
        598 => "00010000",
        599 => "00010000",
        600 => "00010000",
        601 => "00010000",
        602 => "00010000",
        603 => "00010000",
        604 => "00010000",
        605 => "00010000",
        606 => "00010000",
        607 => "00010000",
        608 => "00010000",
        609 => "00010000",
        610 => "00010000",
        611 => "00010000",
        612 => "00010000",
        613 => "00010000",
        614 => "00010000",
        615 => "00010000",
        616 => "00010000",
        617 => "00010000",
        618 => "11011111",
        619 => "11111111",
        620 => "00000001",
        621 => "00000000",
        622 => "11011111",
        623 => "11011111",
        624 => "00110000",
        625 => "00010000",
        626 => "00010000",
        627 => "00010000",
        628 => "00010000",
        629 => "00010000",
        630 => "00010000",
        631 => "00010000",
        632 => "00010000",
        633 => "00010000",
        634 => "00010000",
        635 => "00010000",
        636 => "00010000",
        637 => "00010000",
        638 => "00010000",
        639 => "00010000",
        640 => "00010000",
        641 => "00010000",
        642 => "00010000",
        643 => "00010000",
        644 => "00110000",
        645 => "11011111",
        646 => "11111111",
        647 => "00000001",
        648 => "00000000",
        649 => "10110111",
        650 => "11011111",
        651 => "10011001",
        652 => "00110000",
        653 => "00001100",
        654 => "00101100",
        655 => "00001100",
        656 => "00010000",
        657 => "00010000",
        658 => "00010000",
        659 => "00010000",
        660 => "00010000",
        661 => "00010000",
        662 => "00001100",
        663 => "00001100",
        664 => "00001100",
        665 => "00001100",
        666 => "00010000",
        667 => "00001100",
        668 => "00010000",
        669 => "00001100",
        670 => "00110000",
        671 => "10011010",
        672 => "11011111",
        673 => "10010011",
        674 => "00000001",
        675 => "00000001",
        676 => "00000001",
        677 => "11011111",
        678 => "11011111",
        679 => "11011111",
        680 => "11011111",
        681 => "11011111",
        682 => "11011111",
        683 => "11011111",
        684 => "11011111",
        685 => "11011111",
        686 => "11011111",
        687 => "11011111",
        688 => "11011111",
        689 => "11011111",
        690 => "11011111",
        691 => "11011111",
        692 => "10111111",
        693 => "11011111",
        694 => "11011111",
        695 => "11011111",
        696 => "11011111",
        697 => "11011111",
        698 => "11011111",
        699 => "11011111",
        700 => "00100101",
        701 => "00000001",
        702 => "00000001",
        703 => "00000001",
        704 => "00000101",
        705 => "10010111",
        706 => "11011111",
        707 => "11011111",
        708 => "11111111",
        709 => "11011111",
        710 => "11011111",
        711 => "11011111",
        712 => "11011111",
        713 => "11011111",
        714 => "11011111",
        715 => "11111111",
        716 => "11111111",
        717 => "11111111",
        718 => "11111111",
        719 => "11111111",
        720 => "11111111",
        721 => "11111111",
        722 => "11011111",
        723 => "11011111",
        724 => "11011111",
        725 => "10010111",
        726 => "00100101",
        727 => "00000001",
        728 => "00000001",
        729 => "00000001",
        730 => "00000001",
        731 => "00000001",
        732 => "00000001",
        733 => "00000000",
        734 => "00000000",
        735 => "00000000",
        736 => "00000000",
        737 => "00000000",
        738 => "00000000",
        739 => "00000000",
        740 => "00000000",
        741 => "00000000",
        742 => "00000000",
        743 => "00000000",
        744 => "00000000",
        745 => "00000000",
        746 => "00000000",
        747 => "00000000",
        748 => "00000000",
        749 => "00000000",
        750 => "00000000",
        751 => "00000000",
        752 => "00000000",
        753 => "00000001",
        754 => "00000001",
        755 => "00000001");
        
begin

    process(clk)
    begin
    
        if rising_edge(clk) then
            if rst = '1' then
                Two <= (others => (others => '0'));
            else
                dout <= Two(to_integer(unsigned(addr)));
            end if;
        end if;
    end process;

end Behavioral;



library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity GreenClass is
    port(clk: in std_logic;
         addr: in std_logic_vector(11 downto 0);
         dout: out std_logic_vector(7 downto 0));
end GreenClass;

architecture Behavioral of GreenClass is

    type mem is array (0 to 2623) of std_logic_vector(7 downto 0);
    signal green: mem := (
0 => "00000001",
1 => "00000001",
2 => "00000000",
3 => "00000000",
4 => "00000000",
5 => "00000000",
6 => "00000000",
7 => "00000000",
8 => "00000000",
9 => "00000000",
10 => "00000000",
11 => "00000000",
12 => "00000000",
13 => "00000000",
14 => "00000000",
15 => "00000000",
16 => "00000000",
17 => "00000000",
18 => "00000000",
19 => "00000000",
20 => "00000000",
21 => "00000000",
22 => "00000000",
23 => "00000000",
24 => "00000000",
25 => "00000000",
26 => "00000000",
27 => "00000000",
28 => "00000000",
29 => "00000000",
30 => "00000000",
31 => "00000000",
32 => "00000000",
33 => "00000000",
34 => "00000000",
35 => "00000000",
36 => "00000000",
37 => "00000000",
38 => "00000000",
39 => "00000000",
40 => "00000000",
41 => "00000000",
42 => "00000000",
43 => "00000000",
44 => "00000000",
45 => "00000000",
46 => "00000000",
47 => "00000000",
48 => "00000000",
49 => "00000000",
50 => "00000000",
51 => "00000000",
52 => "00000000",
53 => "00000000",
54 => "00000000",
55 => "00000000",
56 => "00000000",
57 => "00000000",
58 => "00000000",
59 => "00000000",
60 => "00000000",
61 => "00000000",
62 => "00000000",
63 => "00000000",
64 => "00000000",
65 => "00000000",
66 => "00000000",
67 => "00000000",
68 => "00000000",
69 => "00000000",
70 => "00000000",
71 => "00000000",
72 => "00000000",
73 => "00000000",
74 => "00000000",
75 => "00000000",
76 => "00000000",
77 => "00000000",
78 => "00000001",
79 => "00000001",
80 => "00000001",
81 => "00000001",
82 => "00000001",
83 => "00000001",
84 => "00100101",
85 => "10010110",
86 => "11011111",
87 => "11011111",
88 => "11011111",
89 => "11011111",
90 => "11011111",
91 => "11011111",
92 => "11011111",
93 => "11011111",
94 => "11011111",
95 => "11011111",
96 => "11011111",
97 => "11011111",
98 => "11011111",
99 => "11011111",
100 => "11011111",
101 => "11011111",
102 => "11011111",
103 => "11011111",
104 => "11011111",
105 => "11011111",
106 => "11011111",
107 => "11011111",
108 => "11011111",
109 => "11011111",
110 => "11011111",
111 => "11011111",
112 => "11011111",
113 => "11011111",
114 => "11011111",
115 => "11011111",
116 => "11011111",
117 => "11011111",
118 => "11011111",
119 => "11011111",
120 => "11011111",
121 => "11011111",
122 => "11011111",
123 => "11011111",
124 => "11011111",
125 => "11011111",
126 => "11011111",
127 => "11011111",
128 => "11011111",
129 => "11011111",
130 => "11011111",
131 => "11011111",
132 => "11011111",
133 => "11011111",
134 => "11011111",
135 => "11011111",
136 => "11011111",
137 => "11011111",
138 => "11011111",
139 => "11011111",
140 => "11011111",
141 => "11011111",
142 => "11011111",
143 => "11011111",
144 => "11011111",
145 => "11011111",
146 => "11011111",
147 => "11011111",
148 => "11011111",
149 => "11011111",
150 => "11011111",
151 => "11011111",
152 => "11011111",
153 => "11011111",
154 => "11011111",
155 => "11011111",
156 => "11011111",
157 => "11011111",
158 => "11011111",
159 => "11011111",
160 => "10010110",
161 => "00000101",
162 => "00000000",
163 => "00000001",
164 => "00000001",
165 => "00000101",
166 => "10111111",
167 => "01110101",
168 => "00110000",
169 => "00001100",
170 => "00010000",
171 => "00010000",
172 => "00010000",
173 => "00010000",
174 => "00010000",
175 => "00010000",
176 => "00010000",
177 => "00010000",
178 => "00010000",
179 => "00010000",
180 => "00010000",
181 => "00010000",
182 => "00010000",
183 => "00010000",
184 => "00010000",
185 => "00010000",
186 => "00010000",
187 => "00010000",
188 => "00010000",
189 => "00010000",
190 => "00010000",
191 => "00010000",
192 => "00010000",
193 => "00010000",
194 => "00010000",
195 => "00010000",
196 => "00010000",
197 => "00010000",
198 => "00010000",
199 => "00010000",
200 => "00010000",
201 => "00010000",
202 => "00010000",
203 => "00010000",
204 => "00010000",
205 => "00010000",
206 => "00010000",
207 => "00010000",
208 => "00010000",
209 => "00010000",
210 => "00010000",
211 => "00010000",
212 => "00010000",
213 => "00010000",
214 => "00010000",
215 => "00010000",
216 => "00010000",
217 => "00010000",
218 => "00010000",
219 => "00010000",
220 => "00010000",
221 => "00010000",
222 => "00010000",
223 => "00010000",
224 => "00010000",
225 => "00010000",
226 => "00010000",
227 => "00010000",
228 => "00010000",
229 => "00010000",
230 => "00010000",
231 => "00010000",
232 => "00010000",
233 => "00010000",
234 => "00010000",
235 => "00010000",
236 => "00010000",
237 => "00010000",
238 => "00001100",
239 => "00010000",
240 => "00001100",
241 => "00010000",
242 => "01010101",
243 => "10111111",
244 => "00000101",
245 => "00000001",
246 => "00000000",
247 => "10010110",
248 => "01110101",
249 => "00010000",
250 => "00010000",
251 => "00010000",
252 => "00010100",
253 => "00010000",
254 => "00010000",
255 => "00010000",
256 => "00010100",
257 => "00010000",
258 => "00010000",
259 => "00010000",
260 => "00010000",
261 => "00010000",
262 => "00010000",
263 => "00010000",
264 => "00010000",
265 => "00010000",
266 => "00010000",
267 => "00010000",
268 => "00010000",
269 => "00010000",
270 => "00010000",
271 => "00010000",
272 => "00010000",
273 => "00010000",
274 => "00010000",
275 => "00010000",
276 => "00010000",
277 => "00010000",
278 => "00010000",
279 => "00010000",
280 => "00010000",
281 => "00010000",
282 => "00010000",
283 => "00010000",
284 => "00010000",
285 => "00010000",
286 => "00010000",
287 => "00010000",
288 => "00010000",
289 => "00010000",
290 => "00010000",
291 => "00010000",
292 => "00010000",
293 => "00010000",
294 => "00010000",
295 => "00010000",
296 => "00010000",
297 => "00010000",
298 => "00010000",
299 => "00010000",
300 => "00010000",
301 => "00010000",
302 => "00010000",
303 => "00010000",
304 => "00010000",
305 => "00010000",
306 => "00010000",
307 => "00010000",
308 => "00010000",
309 => "00010000",
310 => "00010000",
311 => "00010000",
312 => "00010000",
313 => "00010000",
314 => "00010000",
315 => "00010000",
316 => "00010000",
317 => "00010000",
318 => "00010000",
319 => "00010000",
320 => "00010000",
321 => "00010000",
322 => "00010000",
323 => "00010000",
324 => "00010000",
325 => "01010101",
326 => "10010110",
327 => "00000001",
328 => "00000000",
329 => "11011111",
330 => "00010000",
331 => "00010000",
332 => "00010000",
333 => "00010000",
334 => "00010100",
335 => "00010100",
336 => "00010000",
337 => "00010000",
338 => "00010000",
339 => "00010000",
340 => "00010000",
341 => "00010000",
342 => "00010000",
343 => "00010000",
344 => "00010000",
345 => "00010000",
346 => "00010000",
347 => "00010000",
348 => "00010000",
349 => "00010000",
350 => "00010000",
351 => "00010000",
352 => "00010000",
353 => "00010000",
354 => "00010100",
355 => "00010100",
356 => "00010000",
357 => "00010000",
358 => "00010000",
359 => "00010000",
360 => "00010000",
361 => "00010000",
362 => "00010000",
363 => "00010000",
364 => "00010000",
365 => "00010000",
366 => "00010000",
367 => "00010000",
368 => "00010000",
369 => "00010000",
370 => "00010000",
371 => "00010000",
372 => "00010000",
373 => "00010000",
374 => "00010000",
375 => "00010000",
376 => "00010000",
377 => "00010000",
378 => "00010000",
379 => "00010000",
380 => "00010000",
381 => "00010000",
382 => "00010100",
383 => "00010100",
384 => "00010000",
385 => "00010000",
386 => "00010000",
387 => "00010000",
388 => "00010000",
389 => "00010000",
390 => "00010000",
391 => "00010000",
392 => "00010000",
393 => "00010000",
394 => "00010000",
395 => "00010000",
396 => "00010000",
397 => "00010000",
398 => "00010000",
399 => "00010000",
400 => "00010100",
401 => "00010000",
402 => "00010000",
403 => "00010000",
404 => "00010000",
405 => "00010000",
406 => "00010000",
407 => "00010000",
408 => "11011111",
409 => "00000001",
410 => "00000000",
411 => "11011111",
412 => "00001100",
413 => "00010000",
414 => "00010100",
415 => "00010000",
416 => "00010100",
417 => "00010000",
418 => "00010000",
419 => "00010000",
420 => "00010000",
421 => "00010000",
422 => "00010000",
423 => "00010000",
424 => "00010000",
425 => "00010000",
426 => "00010000",
427 => "00010000",
428 => "00010000",
429 => "00010000",
430 => "00010000",
431 => "00010000",
432 => "00010000",
433 => "00010000",
434 => "00010000",
435 => "00010000",
436 => "00010000",
437 => "00010000",
438 => "00010000",
439 => "00010000",
440 => "00010000",
441 => "00010000",
442 => "00010000",
443 => "00010000",
444 => "00010000",
445 => "00010000",
446 => "00010000",
447 => "00010000",
448 => "00010000",
449 => "00010000",
450 => "00010000",
451 => "00010000",
452 => "00010000",
453 => "00010000",
454 => "00010000",
455 => "00010000",
456 => "00010000",
457 => "00010000",
458 => "00010000",
459 => "00010000",
460 => "00010000",
461 => "00010000",
462 => "00010000",
463 => "00010000",
464 => "00010000",
465 => "00010100",
466 => "00010000",
467 => "00010000",
468 => "00010000",
469 => "00010000",
470 => "00010000",
471 => "00010000",
472 => "00010000",
473 => "00010000",
474 => "00010000",
475 => "00010000",
476 => "00010000",
477 => "00010000",
478 => "00010000",
479 => "00010000",
480 => "00010000",
481 => "00010000",
482 => "00010000",
483 => "00010000",
484 => "00010000",
485 => "00010000",
486 => "00010000",
487 => "00010000",
488 => "00010000",
489 => "00010000",
490 => "11011111",
491 => "00000000",
492 => "00000000",
493 => "11011111",
494 => "00010000",
495 => "00010000",
496 => "00010100",
497 => "00010100",
498 => "00010000",
499 => "00010000",
500 => "00010000",
501 => "00010000",
502 => "00010000",
503 => "00010000",
504 => "00010000",
505 => "00010000",
506 => "00010000",
507 => "00010000",
508 => "00010000",
509 => "00010000",
510 => "00010000",
511 => "00010000",
512 => "00010000",
513 => "00010000",
514 => "00010000",
515 => "00010000",
516 => "00010000",
517 => "00010000",
518 => "00010000",
519 => "00010000",
520 => "00010000",
521 => "00010000",
522 => "00010000",
523 => "00010000",
524 => "00010000",
525 => "00010000",
526 => "00010000",
527 => "00010000",
528 => "00010000",
529 => "00010000",
530 => "00010000",
531 => "00010000",
532 => "00010000",
533 => "00010000",
534 => "00010000",
535 => "00010000",
536 => "00010000",
537 => "00010000",
538 => "00010000",
539 => "00010000",
540 => "00010000",
541 => "00010000",
542 => "00010000",
543 => "00010000",
544 => "00010000",
545 => "00010000",
546 => "00010000",
547 => "00010000",
548 => "00010000",
549 => "00010000",
550 => "00010000",
551 => "00010000",
552 => "00010000",
553 => "00010000",
554 => "00010000",
555 => "00010000",
556 => "00010000",
557 => "00010000",
558 => "00010000",
559 => "00010000",
560 => "00010000",
561 => "00010000",
562 => "00010000",
563 => "00010000",
564 => "00010000",
565 => "00010100",
566 => "00010000",
567 => "00010000",
568 => "00010100",
569 => "00010000",
570 => "00010000",
571 => "00010000",
572 => "11011111",
573 => "00000000",
574 => "00000000",
575 => "11011111",
576 => "00010000",
577 => "00010100",
578 => "00010000",
579 => "00010000",
580 => "00010000",
581 => "00010000",
582 => "00010000",
583 => "00010000",
584 => "00010000",
585 => "00010000",
586 => "00010000",
587 => "00010000",
588 => "00010000",
589 => "00010000",
590 => "00010000",
591 => "00010000",
592 => "00010000",
593 => "00010000",
594 => "00010000",
595 => "00010000",
596 => "00010000",
597 => "00010000",
598 => "00010000",
599 => "00010000",
600 => "00010000",
601 => "00010000",
602 => "00010000",
603 => "00010000",
604 => "00010000",
605 => "00010000",
606 => "00010000",
607 => "00010000",
608 => "00010000",
609 => "00010000",
610 => "00010000",
611 => "00010000",
612 => "00010000",
613 => "00010000",
614 => "00010000",
615 => "00010000",
616 => "00010000",
617 => "00010000",
618 => "00010000",
619 => "00010000",
620 => "00010000",
621 => "00010000",
622 => "00010000",
623 => "00010000",
624 => "00010000",
625 => "00010000",
626 => "00010000",
627 => "00010000",
628 => "00010000",
629 => "00010000",
630 => "00010000",
631 => "00010000",
632 => "00010000",
633 => "00010000",
634 => "00010000",
635 => "00010000",
636 => "00010000",
637 => "00010000",
638 => "00010000",
639 => "00010000",
640 => "00010000",
641 => "00010000",
642 => "00010000",
643 => "00010000",
644 => "00010000",
645 => "00010000",
646 => "00010000",
647 => "00010000",
648 => "00010000",
649 => "00010100",
650 => "00010000",
651 => "00010000",
652 => "00010100",
653 => "00010000",
654 => "11011111",
655 => "00000000",
656 => "00000000",
657 => "11011111",
658 => "00010000",
659 => "00010000",
660 => "00010000",
661 => "00010000",
662 => "00010000",
663 => "00010000",
664 => "00010000",
665 => "00010000",
666 => "00010000",
667 => "00010000",
668 => "00010000",
669 => "00010000",
670 => "00010000",
671 => "00010000",
672 => "00010000",
673 => "00010000",
674 => "00010000",
675 => "00010000",
676 => "00010000",
677 => "00010000",
678 => "00010000",
679 => "00010000",
680 => "00010000",
681 => "00010000",
682 => "00010000",
683 => "00010000",
684 => "00010000",
685 => "00010000",
686 => "00010000",
687 => "00010000",
688 => "00010000",
689 => "00010000",
690 => "00010000",
691 => "00010000",
692 => "00010000",
693 => "00010000",
694 => "00010000",
695 => "00010000",
696 => "00010000",
697 => "00010000",
698 => "00010000",
699 => "00010000",
700 => "00010100",
701 => "00010000",
702 => "00010000",
703 => "00010000",
704 => "00010000",
705 => "00010000",
706 => "00010000",
707 => "00010000",
708 => "00010000",
709 => "00010000",
710 => "00010000",
711 => "00010000",
712 => "00010000",
713 => "00010000",
714 => "00010000",
715 => "00010000",
716 => "00010000",
717 => "00010000",
718 => "00010100",
719 => "00010000",
720 => "00010000",
721 => "00010000",
722 => "00010000",
723 => "00010000",
724 => "00010000",
725 => "00010000",
726 => "00010000",
727 => "00010000",
728 => "00010000",
729 => "00010000",
730 => "00010000",
731 => "00010000",
732 => "00010000",
733 => "00010000",
734 => "00010000",
735 => "00010000",
736 => "11011111",
737 => "00000000",
738 => "00000000",
739 => "11011111",
740 => "00010000",
741 => "00010000",
742 => "00010000",
743 => "00010000",
744 => "00010000",
745 => "00010000",
746 => "00010000",
747 => "00010000",
748 => "00010000",
749 => "00010000",
750 => "00010000",
751 => "00010000",
752 => "00010000",
753 => "00010000",
754 => "00010000",
755 => "00010000",
756 => "00010000",
757 => "00010000",
758 => "00010000",
759 => "00010000",
760 => "00010000",
761 => "00010000",
762 => "00010000",
763 => "00010100",
764 => "00010000",
765 => "00010000",
766 => "00010000",
767 => "00010000",
768 => "00010000",
769 => "00010000",
770 => "00010000",
771 => "00010100",
772 => "00010000",
773 => "00010000",
774 => "00010000",
775 => "00010000",
776 => "00010000",
777 => "00010100",
778 => "00010000",
779 => "00010000",
780 => "00010000",
781 => "00010000",
782 => "00010000",
783 => "00010000",
784 => "00010000",
785 => "00010000",
786 => "00010000",
787 => "00010000",
788 => "00010000",
789 => "00010000",
790 => "00010000",
791 => "00010000",
792 => "00010000",
793 => "00010000",
794 => "00010000",
795 => "00010000",
796 => "00010000",
797 => "00010000",
798 => "00010000",
799 => "00010100",
800 => "00010000",
801 => "00010000",
802 => "00010000",
803 => "00010000",
804 => "00010000",
805 => "00010000",
806 => "00010000",
807 => "00010000",
808 => "00010000",
809 => "00010000",
810 => "00010000",
811 => "00010000",
812 => "00010000",
813 => "00010000",
814 => "00010000",
815 => "00010000",
816 => "00010000",
817 => "00010000",
818 => "11011111",
819 => "00000000",
820 => "00000000",
821 => "11011111",
822 => "00010000",
823 => "00010100",
824 => "00010000",
825 => "00010000",
826 => "00010000",
827 => "00010000",
828 => "00010000",
829 => "00010000",
830 => "00010000",
831 => "00010000",
832 => "00010000",
833 => "00010000",
834 => "00010000",
835 => "00010000",
836 => "00010000",
837 => "00010000",
838 => "00010000",
839 => "00010000",
840 => "00010000",
841 => "00010100",
842 => "00010000",
843 => "00010000",
844 => "00010000",
845 => "00010000",
846 => "00010100",
847 => "00010000",
848 => "00010000",
849 => "00010000",
850 => "00010000",
851 => "00010000",
852 => "00010000",
853 => "00010000",
854 => "00010000",
855 => "00010000",
856 => "00010000",
857 => "00010000",
858 => "00010000",
859 => "00010000",
860 => "00010000",
861 => "00010000",
862 => "00010000",
863 => "00010100",
864 => "00010000",
865 => "00010100",
866 => "00010000",
867 => "00010000",
868 => "00010000",
869 => "00010000",
870 => "00010000",
871 => "00010000",
872 => "00010100",
873 => "00010000",
874 => "00010100",
875 => "00010000",
876 => "00010000",
877 => "00010000",
878 => "00010000",
879 => "00010100",
880 => "00010000",
881 => "00010000",
882 => "00010000",
883 => "00010000",
884 => "00010000",
885 => "00010000",
886 => "00010000",
887 => "00010000",
888 => "00010000",
889 => "00010000",
890 => "00010000",
891 => "00010000",
892 => "00010000",
893 => "00010000",
894 => "00010000",
895 => "00010000",
896 => "00010000",
897 => "00010000",
898 => "00010000",
899 => "00010000",
900 => "11011111",
901 => "00000000",
902 => "00000000",
903 => "11011111",
904 => "00010000",
905 => "00010100",
906 => "00010000",
907 => "00010000",
908 => "00010000",
909 => "00010000",
910 => "00010000",
911 => "00010000",
912 => "00010000",
913 => "00010000",
914 => "00010000",
915 => "00010000",
916 => "00010000",
917 => "00010000",
918 => "00010000",
919 => "00010000",
920 => "00010000",
921 => "00010000",
922 => "00010000",
923 => "00010000",
924 => "00010000",
925 => "00010000",
926 => "00010000",
927 => "00010000",
928 => "00010000",
929 => "00010000",
930 => "00010000",
931 => "00010000",
932 => "00010000",
933 => "00010100",
934 => "00010000",
935 => "00010000",
936 => "00010000",
937 => "00010000",
938 => "00010000",
939 => "00010000",
940 => "00010000",
941 => "00010000",
942 => "00010000",
943 => "00010000",
944 => "00010000",
945 => "00010000",
946 => "00010000",
947 => "00010000",
948 => "00010000",
949 => "00010000",
950 => "00010000",
951 => "00010000",
952 => "00010000",
953 => "00010000",
954 => "00010000",
955 => "00010000",
956 => "00010000",
957 => "00010000",
958 => "00010000",
959 => "00010000",
960 => "00010000",
961 => "00010000",
962 => "00010000",
963 => "00010100",
964 => "00010000",
965 => "00010000",
966 => "00010000",
967 => "00010000",
968 => "00010000",
969 => "00010000",
970 => "00010000",
971 => "00010000",
972 => "00010000",
973 => "00010000",
974 => "00010000",
975 => "00010000",
976 => "00010000",
977 => "00010000",
978 => "00010000",
979 => "00010000",
980 => "00010000",
981 => "00010000",
982 => "11011111",
983 => "00000000",
984 => "00000000",
985 => "11011111",
986 => "00010000",
987 => "00010000",
988 => "00010000",
989 => "00010000",
990 => "00010000",
991 => "00010000",
992 => "00010000",
993 => "00010000",
994 => "00010000",
995 => "00010000",
996 => "00010000",
997 => "00010000",
998 => "00010000",
999 => "00010000",
1000 => "00010000",
1001 => "00010000",
1002 => "00010000",
1003 => "00010000",
1004 => "00010000",
1005 => "00010100",
1006 => "10111110",
1007 => "11011110",
1008 => "01010100",
1009 => "00001100",
1010 => "10011110",
1011 => "10011110",
1012 => "00010000",
1013 => "00010100",
1014 => "00010000",
1015 => "00010000",
1016 => "00010000",
1017 => "00010000",
1018 => "00010000",
1019 => "00010100",
1020 => "00010000",
1021 => "00010000",
1022 => "00010000",
1023 => "00010000",
1024 => "00010000",
1025 => "00010000",
1026 => "00010000",
1027 => "00010000",
1028 => "00010000",
1029 => "00010000",
1030 => "00010000",
1031 => "00010000",
1032 => "00010000",
1033 => "00010000",
1034 => "00010000",
1035 => "00010000",
1036 => "00010000",
1037 => "00010000",
1038 => "00010000",
1039 => "01011101",
1040 => "10111110",
1041 => "11011110",
1042 => "10111110",
1043 => "01010100",
1044 => "00010000",
1045 => "00010000",
1046 => "00010000",
1047 => "00010000",
1048 => "00010000",
1049 => "00010000",
1050 => "00010000",
1051 => "00010000",
1052 => "00010000",
1053 => "00010000",
1054 => "00010000",
1055 => "00010000",
1056 => "00010000",
1057 => "00010000",
1058 => "00010000",
1059 => "00010000",
1060 => "00010000",
1061 => "00010000",
1062 => "00010000",
1063 => "00010000",
1064 => "11011111",
1065 => "00000000",
1066 => "00000000",
1067 => "11011111",
1068 => "00010000",
1069 => "00010000",
1070 => "00010000",
1071 => "00010000",
1072 => "00010000",
1073 => "00010000",
1074 => "00010000",
1075 => "00010000",
1076 => "00010000",
1077 => "00010000",
1078 => "00010000",
1079 => "00010000",
1080 => "00010000",
1081 => "00010000",
1082 => "00010000",
1083 => "00010000",
1084 => "00010000",
1085 => "00010000",
1086 => "00010000",
1087 => "00010000",
1088 => "11011111",
1089 => "11111111",
1090 => "10111101",
1091 => "01001100",
1092 => "10111110",
1093 => "10111110",
1094 => "00010000",
1095 => "00010000",
1096 => "00010000",
1097 => "00010000",
1098 => "00010000",
1099 => "00010000",
1100 => "00010000",
1101 => "00010000",
1102 => "00010000",
1103 => "00010000",
1104 => "00010000",
1105 => "00010000",
1106 => "00010000",
1107 => "00010000",
1108 => "00010000",
1109 => "00010000",
1110 => "00010000",
1111 => "00010000",
1112 => "00010000",
1113 => "00010000",
1114 => "00010000",
1115 => "00010000",
1116 => "00010000",
1117 => "00010000",
1118 => "00010000",
1119 => "00010000",
1120 => "00010000",
1121 => "00010000",
1122 => "00110000",
1123 => "10111110",
1124 => "11011110",
1125 => "01010000",
1126 => "00010000",
1127 => "00010000",
1128 => "00010100",
1129 => "00010000",
1130 => "00010000",
1131 => "00010000",
1132 => "00010000",
1133 => "00010000",
1134 => "00010000",
1135 => "00010000",
1136 => "00010000",
1137 => "00010000",
1138 => "00010000",
1139 => "00010000",
1140 => "00010000",
1141 => "00010000",
1142 => "00010000",
1143 => "00010000",
1144 => "00010000",
1145 => "00010000",
1146 => "11011111",
1147 => "00000000",
1148 => "00000000",
1149 => "11011111",
1150 => "00010000",
1151 => "00010000",
1152 => "00010000",
1153 => "00010000",
1154 => "00010000",
1155 => "00010000",
1156 => "00010000",
1157 => "00010000",
1158 => "00010000",
1159 => "00010000",
1160 => "00010000",
1161 => "00010000",
1162 => "00010000",
1163 => "00010000",
1164 => "00010000",
1165 => "00010000",
1166 => "00010000",
1167 => "00010000",
1168 => "00010000",
1169 => "00010000",
1170 => "10111111",
1171 => "11011110",
1172 => "11111110",
1173 => "10010000",
1174 => "10111010",
1175 => "10111110",
1176 => "00010000",
1177 => "00010000",
1178 => "10111110",
1179 => "11011110",
1180 => "11011110",
1181 => "10011110",
1182 => "00010000",
1183 => "00110101",
1184 => "10111110",
1185 => "10111110",
1186 => "11011110",
1187 => "10111110",
1188 => "10011110",
1189 => "01010101",
1190 => "11011110",
1191 => "11011110",
1192 => "11011110",
1193 => "10111110",
1194 => "11011110",
1195 => "10111110",
1196 => "00010000",
1197 => "10011110",
1198 => "10111110",
1199 => "10111110",
1200 => "11011110",
1201 => "01111001",
1202 => "00010000",
1203 => "00010000",
1204 => "00110001",
1205 => "10111110",
1206 => "11011110",
1207 => "01010000",
1208 => "00010000",
1209 => "00010000",
1210 => "00010000",
1211 => "00010000",
1212 => "00010000",
1213 => "00010000",
1214 => "00010000",
1215 => "00010000",
1216 => "00010000",
1217 => "00010000",
1218 => "00010000",
1219 => "00010000",
1220 => "00010000",
1221 => "00010000",
1222 => "00010000",
1223 => "00010000",
1224 => "00010000",
1225 => "00010000",
1226 => "00010000",
1227 => "00010000",
1228 => "11011111",
1229 => "00000000",
1230 => "00000000",
1231 => "11011111",
1232 => "00010000",
1233 => "00010000",
1234 => "00010000",
1235 => "00010000",
1236 => "00010000",
1237 => "00010000",
1238 => "00010000",
1239 => "00010000",
1240 => "00010000",
1241 => "00010000",
1242 => "00010000",
1243 => "00010000",
1244 => "00010000",
1245 => "00010000",
1246 => "00010000",
1247 => "00010000",
1248 => "00010000",
1249 => "00010000",
1250 => "00010000",
1251 => "00010000",
1252 => "10111110",
1253 => "11011110",
1254 => "11111110",
1255 => "10110101",
1256 => "10111010",
1257 => "10111110",
1258 => "00010001",
1259 => "10011110",
1260 => "10111110",
1261 => "00101100",
1262 => "01110101",
1263 => "10111111",
1264 => "01111110",
1265 => "00110101",
1266 => "11011110",
1267 => "11011110",
1268 => "01010000",
1269 => "01111001",
1270 => "10111110",
1271 => "01111010",
1272 => "11011110",
1273 => "11011010",
1274 => "11011110",
1275 => "11011110",
1276 => "10111010",
1277 => "10111110",
1278 => "00001100",
1279 => "00001100",
1280 => "00101100",
1281 => "00101100",
1282 => "10111010",
1283 => "11011110",
1284 => "00110100",
1285 => "00010000",
1286 => "00010001",
1287 => "10111111",
1288 => "11011110",
1289 => "01010100",
1290 => "00010000",
1291 => "00010000",
1292 => "00010000",
1293 => "00010000",
1294 => "00010000",
1295 => "00010000",
1296 => "00010000",
1297 => "00010000",
1298 => "00010000",
1299 => "00010000",
1300 => "00010000",
1301 => "00010000",
1302 => "00010000",
1303 => "00010000",
1304 => "00010000",
1305 => "00010000",
1306 => "00010000",
1307 => "00010000",
1308 => "00010000",
1309 => "00010000",
1310 => "11011111",
1311 => "00000000",
1312 => "00000000",
1313 => "11011111",
1314 => "00010000",
1315 => "00010000",
1316 => "00010000",
1317 => "00010000",
1318 => "00010000",
1319 => "00010000",
1320 => "00010000",
1321 => "00010000",
1322 => "00010000",
1323 => "00010000",
1324 => "00010000",
1325 => "00010000",
1326 => "00010000",
1327 => "00010000",
1328 => "00010000",
1329 => "00010000",
1330 => "00010000",
1331 => "00010000",
1332 => "00010000",
1333 => "00010000",
1334 => "11011110",
1335 => "10111001",
1336 => "10111010",
1337 => "11011111",
1338 => "11011110",
1339 => "10111110",
1340 => "00110101",
1341 => "10111110",
1342 => "10011001",
1343 => "00101100",
1344 => "00110001",
1345 => "10011111",
1346 => "10011110",
1347 => "01010100",
1348 => "11011110",
1349 => "10111001",
1350 => "00010000",
1351 => "00010000",
1352 => "00010000",
1353 => "00110101",
1354 => "11011110",
1355 => "10110101",
1356 => "11011110",
1357 => "10111010",
1358 => "10011010",
1359 => "11011111",
1360 => "01010001",
1361 => "10011001",
1362 => "11011110",
1363 => "11011110",
1364 => "11111110",
1365 => "11011110",
1366 => "01010100",
1367 => "00010000",
1368 => "00110000",
1369 => "10111110",
1370 => "11011110",
1371 => "01010000",
1372 => "00010000",
1373 => "00010000",
1374 => "00010000",
1375 => "00010000",
1376 => "00010000",
1377 => "00010000",
1378 => "00010000",
1379 => "00010000",
1380 => "00010000",
1381 => "00010000",
1382 => "00010000",
1383 => "00010000",
1384 => "00010000",
1385 => "00010000",
1386 => "00010000",
1387 => "00010000",
1388 => "00010000",
1389 => "00010000",
1390 => "00010000",
1391 => "00010000",
1392 => "11011111",
1393 => "00000000",
1394 => "00000000",
1395 => "11011111",
1396 => "00010000",
1397 => "00010000",
1398 => "00010000",
1399 => "00010000",
1400 => "00010000",
1401 => "00010000",
1402 => "00010000",
1403 => "00010000",
1404 => "00010000",
1405 => "00010000",
1406 => "00010000",
1407 => "00010000",
1408 => "00010000",
1409 => "00010000",
1410 => "00010000",
1411 => "00010000",
1412 => "00010100",
1413 => "00010000",
1414 => "00010000",
1415 => "00010000",
1416 => "11011110",
1417 => "10111001",
1418 => "01010001",
1419 => "10111111",
1420 => "11011111",
1421 => "11011110",
1422 => "00110101",
1423 => "10011111",
1424 => "10011001",
1425 => "00101100",
1426 => "00101100",
1427 => "10111111",
1428 => "10011110",
1429 => "01010101",
1430 => "11011101",
1431 => "10011000",
1432 => "00010000",
1433 => "00010000",
1434 => "00010000",
1435 => "00110101",
1436 => "11011110",
1437 => "10110101",
1438 => "11011110",
1439 => "10111010",
1440 => "10011010",
1441 => "10111111",
1442 => "10011010",
1443 => "11011110",
1444 => "10011001",
1445 => "00101100",
1446 => "10111010",
1447 => "11011110",
1448 => "01010000",
1449 => "00010000",
1450 => "00110000",
1451 => "10111110",
1452 => "11011110",
1453 => "01010000",
1454 => "00010000",
1455 => "00010000",
1456 => "00010000",
1457 => "00010000",
1458 => "00010000",
1459 => "00010000",
1460 => "00010000",
1461 => "00010000",
1462 => "00010000",
1463 => "00010000",
1464 => "00010000",
1465 => "00010000",
1466 => "00010000",
1467 => "00010000",
1468 => "00010000",
1469 => "00010000",
1470 => "00010000",
1471 => "00010000",
1472 => "00010000",
1473 => "00010000",
1474 => "11011111",
1475 => "00000000",
1476 => "00000000",
1477 => "11011111",
1478 => "00010000",
1479 => "00010000",
1480 => "00010000",
1481 => "00010000",
1482 => "00010000",
1483 => "00010000",
1484 => "00010000",
1485 => "00010000",
1486 => "00010000",
1487 => "00010000",
1488 => "00010000",
1489 => "00010000",
1490 => "00010000",
1491 => "00010000",
1492 => "00010000",
1493 => "00010000",
1494 => "00010000",
1495 => "00010000",
1496 => "00010000",
1497 => "00010000",
1498 => "11011110",
1499 => "10011001",
1500 => "00010000",
1501 => "10011111",
1502 => "11011111",
1503 => "11011110",
1504 => "00010001",
1505 => "10011110",
1506 => "10111110",
1507 => "00101100",
1508 => "01110101",
1509 => "10111111",
1510 => "01011001",
1511 => "01010100",
1512 => "11111110",
1513 => "10111001",
1514 => "00010000",
1515 => "00010000",
1516 => "00010000",
1517 => "00110101",
1518 => "11011110",
1519 => "10110101",
1520 => "11011110",
1521 => "10111110",
1522 => "10011010",
1523 => "11011111",
1524 => "10011010",
1525 => "11011111",
1526 => "01110101",
1527 => "01110001",
1528 => "11011111",
1529 => "11011110",
1530 => "01010000",
1531 => "00101100",
1532 => "00110000",
1533 => "10111110",
1534 => "11011110",
1535 => "01010000",
1536 => "00010000",
1537 => "00010000",
1538 => "00010000",
1539 => "00010000",
1540 => "00010000",
1541 => "00010000",
1542 => "00010000",
1543 => "00010000",
1544 => "00010000",
1545 => "00010000",
1546 => "00010000",
1547 => "00010000",
1548 => "00010000",
1549 => "00010000",
1550 => "00010000",
1551 => "00010000",
1552 => "00010000",
1553 => "00010000",
1554 => "00010000",
1555 => "00010000",
1556 => "11011111",
1557 => "00000000",
1558 => "00000000",
1559 => "11011111",
1560 => "00010000",
1561 => "00010000",
1562 => "00010000",
1563 => "00010000",
1564 => "00010000",
1565 => "00010000",
1566 => "00010000",
1567 => "00010000",
1568 => "00010000",
1569 => "00010000",
1570 => "00010000",
1571 => "00010000",
1572 => "00010000",
1573 => "00010000",
1574 => "00010000",
1575 => "00010000",
1576 => "00010000",
1577 => "00010000",
1578 => "00010000",
1579 => "00010000",
1580 => "10111110",
1581 => "10011001",
1582 => "00010000",
1583 => "00110101",
1584 => "11011110",
1585 => "10111110",
1586 => "00001100",
1587 => "00110101",
1588 => "10111110",
1589 => "10111110",
1590 => "10111110",
1591 => "01111101",
1592 => "00010000",
1593 => "00110100",
1594 => "11011110",
1595 => "10011000",
1596 => "00010000",
1597 => "00010000",
1598 => "00010000",
1599 => "00010100",
1600 => "10111110",
1601 => "10011001",
1602 => "10111101",
1603 => "10111110",
1604 => "10011001",
1605 => "10111110",
1606 => "01010101",
1607 => "10111110",
1608 => "10111110",
1609 => "10111110",
1610 => "10011110",
1611 => "10111110",
1612 => "01010000",
1613 => "10011101",
1614 => "10111110",
1615 => "10111110",
1616 => "10111110",
1617 => "10111110",
1618 => "10011101",
1619 => "00010000",
1620 => "00010000",
1621 => "00010000",
1622 => "00010000",
1623 => "00010000",
1624 => "00010000",
1625 => "00010000",
1626 => "00010000",
1627 => "00010000",
1628 => "00010000",
1629 => "00010000",
1630 => "00010000",
1631 => "00010000",
1632 => "00010000",
1633 => "00010000",
1634 => "00010000",
1635 => "00010000",
1636 => "00010000",
1637 => "00010000",
1638 => "11011111",
1639 => "00000000",
1640 => "00000000",
1641 => "11011111",
1642 => "00010000",
1643 => "00010100",
1644 => "00010000",
1645 => "00010000",
1646 => "00010000",
1647 => "00010000",
1648 => "00010000",
1649 => "00010000",
1650 => "00010000",
1651 => "00010000",
1652 => "00010000",
1653 => "00010000",
1654 => "00010000",
1655 => "00010000",
1656 => "00010000",
1657 => "00010100",
1658 => "00010100",
1659 => "00010000",
1660 => "00010000",
1661 => "00010000",
1662 => "00010000",
1663 => "00010000",
1664 => "00010000",
1665 => "00010000",
1666 => "00010000",
1667 => "00010000",
1668 => "00010000",
1669 => "00010000",
1670 => "00010000",
1671 => "00010000",
1672 => "00010000",
1673 => "00010000",
1674 => "00010000",
1675 => "00010000",
1676 => "00010000",
1677 => "00010000",
1678 => "00010000",
1679 => "00010000",
1680 => "00010000",
1681 => "00010000",
1682 => "00010000",
1683 => "00010000",
1684 => "00010000",
1685 => "00010000",
1686 => "00010000",
1687 => "00010000",
1688 => "00010000",
1689 => "00010000",
1690 => "00010000",
1691 => "00010000",
1692 => "00010000",
1693 => "00010000",
1694 => "00010000",
1695 => "00010000",
1696 => "00010000",
1697 => "00010000",
1698 => "00010000",
1699 => "00010000",
1700 => "00010000",
1701 => "00010100",
1702 => "00010000",
1703 => "00010000",
1704 => "00010000",
1705 => "00010000",
1706 => "00010000",
1707 => "00010000",
1708 => "00010000",
1709 => "00010000",
1710 => "00010000",
1711 => "00010000",
1712 => "00010000",
1713 => "00010000",
1714 => "00010000",
1715 => "00010000",
1716 => "00010000",
1717 => "00010000",
1718 => "00010000",
1719 => "00010000",
1720 => "11011111",
1721 => "00000000",
1722 => "00000000",
1723 => "11011111",
1724 => "00010000",
1725 => "00010100",
1726 => "00010000",
1727 => "00010000",
1728 => "00010000",
1729 => "00010000",
1730 => "00010000",
1731 => "00010000",
1732 => "00010000",
1733 => "00010000",
1734 => "00010000",
1735 => "00010000",
1736 => "00010000",
1737 => "00010000",
1738 => "00010000",
1739 => "00010000",
1740 => "00010000",
1741 => "00010000",
1742 => "00010000",
1743 => "00010000",
1744 => "00010000",
1745 => "00010000",
1746 => "00010000",
1747 => "00010000",
1748 => "00010000",
1749 => "00010000",
1750 => "00010000",
1751 => "00010000",
1752 => "00010000",
1753 => "00010000",
1754 => "00010000",
1755 => "00010000",
1756 => "00010000",
1757 => "00010000",
1758 => "00010000",
1759 => "00010000",
1760 => "00010000",
1761 => "00010000",
1762 => "00010000",
1763 => "00010000",
1764 => "00010100",
1765 => "00010100",
1766 => "00010000",
1767 => "00010000",
1768 => "00010000",
1769 => "00010000",
1770 => "00010000",
1771 => "00010100",
1772 => "00010000",
1773 => "00010000",
1774 => "00010100",
1775 => "00010000",
1776 => "00010000",
1777 => "00010000",
1778 => "00010000",
1779 => "00010000",
1780 => "00010000",
1781 => "00010100",
1782 => "00010000",
1783 => "00010000",
1784 => "00010100",
1785 => "00010000",
1786 => "00010000",
1787 => "00010000",
1788 => "00010000",
1789 => "00010000",
1790 => "00010000",
1791 => "00010000",
1792 => "00010000",
1793 => "00010000",
1794 => "00010000",
1795 => "00010000",
1796 => "00010000",
1797 => "00010000",
1798 => "00010000",
1799 => "00010000",
1800 => "00010000",
1801 => "00010000",
1802 => "11011111",
1803 => "00000000",
1804 => "00000000",
1805 => "11011111",
1806 => "00010000",
1807 => "00010000",
1808 => "00010000",
1809 => "00010000",
1810 => "00010000",
1811 => "00010000",
1812 => "00010000",
1813 => "00010000",
1814 => "00010000",
1815 => "00010000",
1816 => "00010000",
1817 => "00010000",
1818 => "00010000",
1819 => "00010000",
1820 => "00010000",
1821 => "00010000",
1822 => "00010000",
1823 => "00010000",
1824 => "00010000",
1825 => "00010000",
1826 => "00010000",
1827 => "00010000",
1828 => "00010000",
1829 => "00010000",
1830 => "00010000",
1831 => "00010100",
1832 => "00010000",
1833 => "00010000",
1834 => "00010000",
1835 => "00010000",
1836 => "00010000",
1837 => "00010100",
1838 => "00010000",
1839 => "00010000",
1840 => "00010000",
1841 => "00010000",
1842 => "00010000",
1843 => "00010100",
1844 => "00010000",
1845 => "00010000",
1846 => "00010000",
1847 => "00010000",
1848 => "00010000",
1849 => "00010000",
1850 => "00010000",
1851 => "00010000",
1852 => "00010000",
1853 => "00010000",
1854 => "00010100",
1855 => "00010000",
1856 => "00010000",
1857 => "00010000",
1858 => "00010000",
1859 => "00010000",
1860 => "00010000",
1861 => "00010000",
1862 => "00010000",
1863 => "00010000",
1864 => "00010000",
1865 => "00010100",
1866 => "00010000",
1867 => "00010000",
1868 => "00010000",
1869 => "00010000",
1870 => "00010000",
1871 => "00010000",
1872 => "00010000",
1873 => "00010000",
1874 => "00010000",
1875 => "00010000",
1876 => "00010000",
1877 => "00010000",
1878 => "00010000",
1879 => "00010000",
1880 => "00010000",
1881 => "00010000",
1882 => "00010000",
1883 => "00010000",
1884 => "11011111",
1885 => "00000000",
1886 => "00000000",
1887 => "11011111",
1888 => "00010000",
1889 => "00010000",
1890 => "00010000",
1891 => "00010000",
1892 => "00010000",
1893 => "00010000",
1894 => "00010000",
1895 => "00010000",
1896 => "00010000",
1897 => "00010000",
1898 => "00010000",
1899 => "00010000",
1900 => "00010000",
1901 => "00010000",
1902 => "00010000",
1903 => "00010000",
1904 => "00010000",
1905 => "00010000",
1906 => "00010000",
1907 => "00010000",
1908 => "00010000",
1909 => "00010100",
1910 => "00010000",
1911 => "00010100",
1912 => "00010000",
1913 => "00010000",
1914 => "00010000",
1915 => "00010000",
1916 => "00010000",
1917 => "00010000",
1918 => "00010000",
1919 => "00010000",
1920 => "00010000",
1921 => "00010000",
1922 => "00010000",
1923 => "00010000",
1924 => "00010000",
1925 => "00010000",
1926 => "00010000",
1927 => "00010100",
1928 => "00010000",
1929 => "00010000",
1930 => "00010000",
1931 => "00010000",
1932 => "00010000",
1933 => "00010000",
1934 => "00010000",
1935 => "00010000",
1936 => "00010000",
1937 => "00010100",
1938 => "00010000",
1939 => "00010000",
1940 => "00010000",
1941 => "00010000",
1942 => "00010000",
1943 => "00010000",
1944 => "00010000",
1945 => "00010000",
1946 => "00010000",
1947 => "00010000",
1948 => "00010000",
1949 => "00010000",
1950 => "00010000",
1951 => "00010000",
1952 => "00010000",
1953 => "00010000",
1954 => "00010000",
1955 => "00010000",
1956 => "00010000",
1957 => "00010000",
1958 => "00010000",
1959 => "00010000",
1960 => "00010000",
1961 => "00010000",
1962 => "00010000",
1963 => "00010000",
1964 => "00010000",
1965 => "00010000",
1966 => "11011111",
1967 => "00000000",
1968 => "00000000",
1969 => "11011111",
1970 => "00010000",
1971 => "00010100",
1972 => "00010000",
1973 => "00010000",
1974 => "00010000",
1975 => "00010000",
1976 => "00010000",
1977 => "00010000",
1978 => "00010000",
1979 => "00010000",
1980 => "00010000",
1981 => "00010000",
1982 => "00010000",
1983 => "00010000",
1984 => "00010000",
1985 => "00010000",
1986 => "00010000",
1987 => "00010000",
1988 => "00010000",
1989 => "00010000",
1990 => "00010000",
1991 => "00010000",
1992 => "00010000",
1993 => "00010000",
1994 => "00010000",
1995 => "00010000",
1996 => "00010000",
1997 => "00010000",
1998 => "00010000",
1999 => "00010000",
2000 => "00010000",
2001 => "00010000",
2002 => "00010000",
2003 => "00010000",
2004 => "00010000",
2005 => "00010000",
2006 => "00010000",
2007 => "00010000",
2008 => "00010000",
2009 => "00010000",
2010 => "00010000",
2011 => "00010000",
2012 => "00010000",
2013 => "00010000",
2014 => "00010000",
2015 => "00010000",
2016 => "00010000",
2017 => "00010000",
2018 => "00010000",
2019 => "00010000",
2020 => "00010000",
2021 => "00010000",
2022 => "00010000",
2023 => "00010000",
2024 => "00010000",
2025 => "00010000",
2026 => "00010000",
2027 => "00010000",
2028 => "00010000",
2029 => "00010000",
2030 => "00010000",
2031 => "00010000",
2032 => "00010000",
2033 => "00010000",
2034 => "00010000",
2035 => "00010000",
2036 => "00010000",
2037 => "00010000",
2038 => "00010000",
2039 => "00010000",
2040 => "00010000",
2041 => "00010000",
2042 => "00010000",
2043 => "00010100",
2044 => "00010000",
2045 => "00010000",
2046 => "00010100",
2047 => "00010000",
2048 => "11011111",
2049 => "00000000",
2050 => "00000000",
2051 => "11011111",
2052 => "00010000",
2053 => "00010000",
2054 => "00010100",
2055 => "00010100",
2056 => "00010000",
2057 => "00010000",
2058 => "00010000",
2059 => "00010000",
2060 => "00010000",
2061 => "00010000",
2062 => "00010000",
2063 => "00010000",
2064 => "00010000",
2065 => "00010000",
2066 => "00010000",
2067 => "00010000",
2068 => "00010000",
2069 => "00010000",
2070 => "00010000",
2071 => "00010000",
2072 => "00010000",
2073 => "00010000",
2074 => "00010000",
2075 => "00010000",
2076 => "00010000",
2077 => "00010000",
2078 => "00010000",
2079 => "00010000",
2080 => "00010000",
2081 => "00010000",
2082 => "00010000",
2083 => "00010000",
2084 => "00010000",
2085 => "00010000",
2086 => "00010000",
2087 => "00010000",
2088 => "00010000",
2089 => "00010000",
2090 => "00010000",
2091 => "00010000",
2092 => "00010000",
2093 => "00010000",
2094 => "00010000",
2095 => "00010000",
2096 => "00010000",
2097 => "00010000",
2098 => "00010000",
2099 => "00010000",
2100 => "00010000",
2101 => "00010000",
2102 => "00010000",
2103 => "00010000",
2104 => "00010000",
2105 => "00010000",
2106 => "00010000",
2107 => "00010000",
2108 => "00010000",
2109 => "00010000",
2110 => "00010000",
2111 => "00010000",
2112 => "00010000",
2113 => "00010000",
2114 => "00010000",
2115 => "00010000",
2116 => "00010000",
2117 => "00010000",
2118 => "00010000",
2119 => "00010000",
2120 => "00010000",
2121 => "00010000",
2122 => "00010000",
2123 => "00010100",
2124 => "00010000",
2125 => "00010000",
2126 => "00010100",
2127 => "00010000",
2128 => "00010000",
2129 => "00010000",
2130 => "11011111",
2131 => "00000000",
2132 => "00000000",
2133 => "11011111",
2134 => "00001100",
2135 => "00010000",
2136 => "00010100",
2137 => "00010000",
2138 => "00010100",
2139 => "00010000",
2140 => "00010000",
2141 => "00010000",
2142 => "00010000",
2143 => "00010000",
2144 => "00010000",
2145 => "00010000",
2146 => "00010000",
2147 => "00010000",
2148 => "00010000",
2149 => "00010000",
2150 => "00010000",
2151 => "00010000",
2152 => "00010000",
2153 => "00010000",
2154 => "00010000",
2155 => "00010000",
2156 => "00010000",
2157 => "00010000",
2158 => "00010000",
2159 => "00010000",
2160 => "00010000",
2161 => "00010000",
2162 => "00010000",
2163 => "00010000",
2164 => "00010000",
2165 => "00010000",
2166 => "00010000",
2167 => "00010000",
2168 => "00010000",
2169 => "00010000",
2170 => "00010000",
2171 => "00010000",
2172 => "00010000",
2173 => "00010000",
2174 => "00010000",
2175 => "00010000",
2176 => "00010000",
2177 => "00010000",
2178 => "00010000",
2179 => "00010000",
2180 => "00010000",
2181 => "00010000",
2182 => "00010000",
2183 => "00010000",
2184 => "00010000",
2185 => "00010000",
2186 => "00010000",
2187 => "00010000",
2188 => "00010000",
2189 => "00010000",
2190 => "00010000",
2191 => "00010000",
2192 => "00010000",
2193 => "00010000",
2194 => "00010000",
2195 => "00010000",
2196 => "00010000",
2197 => "00010000",
2198 => "00010000",
2199 => "00010000",
2200 => "00010000",
2201 => "00010000",
2202 => "00010000",
2203 => "00010000",
2204 => "00010000",
2205 => "00010000",
2206 => "00010000",
2207 => "00010000",
2208 => "00010000",
2209 => "00010000",
2210 => "00010000",
2211 => "00010000",
2212 => "11011111",
2213 => "00000000",
2214 => "00000000",
2215 => "11011111",
2216 => "00010000",
2217 => "00010000",
2218 => "00010000",
2219 => "00010000",
2220 => "00010100",
2221 => "00010100",
2222 => "00010000",
2223 => "00010000",
2224 => "00010000",
2225 => "00010000",
2226 => "00010000",
2227 => "00010000",
2228 => "00010000",
2229 => "00010000",
2230 => "00010000",
2231 => "00010000",
2232 => "00010000",
2233 => "00010000",
2234 => "00010000",
2235 => "00010000",
2236 => "00010000",
2237 => "00010000",
2238 => "00010000",
2239 => "00010000",
2240 => "00010000",
2241 => "00010000",
2242 => "00010000",
2243 => "00010000",
2244 => "00010100",
2245 => "00010100",
2246 => "00010000",
2247 => "00010000",
2248 => "00010000",
2249 => "00010000",
2250 => "00010000",
2251 => "00010000",
2252 => "00010000",
2253 => "00010000",
2254 => "00010000",
2255 => "00010000",
2256 => "00010000",
2257 => "00010000",
2258 => "00010000",
2259 => "00010000",
2260 => "00010000",
2261 => "00010000",
2262 => "00010000",
2263 => "00010000",
2264 => "00010000",
2265 => "00010000",
2266 => "00010000",
2267 => "00010000",
2268 => "00010000",
2269 => "00010000",
2270 => "00010000",
2271 => "00010000",
2272 => "00010000",
2273 => "00010000",
2274 => "00010000",
2275 => "00010000",
2276 => "00010000",
2277 => "00010000",
2278 => "00010000",
2279 => "00010000",
2280 => "00010000",
2281 => "00010000",
2282 => "00010000",
2283 => "00010000",
2284 => "00010000",
2285 => "00010000",
2286 => "00010100",
2287 => "00010000",
2288 => "00010000",
2289 => "00010000",
2290 => "00010000",
2291 => "00010000",
2292 => "00010000",
2293 => "00010000",
2294 => "11011111",
2295 => "00000001",
2296 => "00000000",
2297 => "10010110",
2298 => "01110101",
2299 => "00010000",
2300 => "00010000",
2301 => "00010000",
2302 => "00010100",
2303 => "00010000",
2304 => "00010000",
2305 => "00010000",
2306 => "00010100",
2307 => "00010000",
2308 => "00010000",
2309 => "00010000",
2310 => "00010000",
2311 => "00010000",
2312 => "00010000",
2313 => "00010000",
2314 => "00010000",
2315 => "00010000",
2316 => "00010000",
2317 => "00010000",
2318 => "00010000",
2319 => "00010000",
2320 => "00010000",
2321 => "00010000",
2322 => "00010000",
2323 => "00010000",
2324 => "00010000",
2325 => "00010000",
2326 => "00010000",
2327 => "00010000",
2328 => "00010000",
2329 => "00010000",
2330 => "00010000",
2331 => "00010000",
2332 => "00010000",
2333 => "00010000",
2334 => "00010000",
2335 => "00010000",
2336 => "00010000",
2337 => "00010000",
2338 => "00010000",
2339 => "00010000",
2340 => "00010000",
2341 => "00010000",
2342 => "00010000",
2343 => "00010000",
2344 => "00010000",
2345 => "00010000",
2346 => "00010000",
2347 => "00010000",
2348 => "00010000",
2349 => "00010000",
2350 => "00010000",
2351 => "00010000",
2352 => "00010000",
2353 => "00010000",
2354 => "00010000",
2355 => "00010000",
2356 => "00010000",
2357 => "00010000",
2358 => "00010000",
2359 => "00010000",
2360 => "00010000",
2361 => "00010000",
2362 => "00010000",
2363 => "00010000",
2364 => "00010000",
2365 => "00010000",
2366 => "00010000",
2367 => "00010000",
2368 => "00010000",
2369 => "00010000",
2370 => "00010000",
2371 => "00010000",
2372 => "00010000",
2373 => "00010000",
2374 => "00010000",
2375 => "01010101",
2376 => "10010110",
2377 => "00000001",
2378 => "00000001",
2379 => "00000101",
2380 => "10111111",
2381 => "01110101",
2382 => "00110000",
2383 => "00001100",
2384 => "00010000",
2385 => "00010000",
2386 => "00010000",
2387 => "00010000",
2388 => "00010000",
2389 => "00010000",
2390 => "00010000",
2391 => "00010000",
2392 => "00010000",
2393 => "00010000",
2394 => "00010000",
2395 => "00010000",
2396 => "00010000",
2397 => "00010000",
2398 => "00010000",
2399 => "00010000",
2400 => "00010000",
2401 => "00010000",
2402 => "00010000",
2403 => "00010000",
2404 => "00010000",
2405 => "00010000",
2406 => "00010000",
2407 => "00010000",
2408 => "00010000",
2409 => "00010000",
2410 => "00010000",
2411 => "00010000",
2412 => "00010000",
2413 => "00010000",
2414 => "00010000",
2415 => "00010000",
2416 => "00010000",
2417 => "00010000",
2418 => "00010000",
2419 => "00010000",
2420 => "00010000",
2421 => "00010000",
2422 => "00010000",
2423 => "00010000",
2424 => "00010000",
2425 => "00010000",
2426 => "00010000",
2427 => "00010000",
2428 => "00010000",
2429 => "00010000",
2430 => "00010000",
2431 => "00010000",
2432 => "00010000",
2433 => "00010000",
2434 => "00010000",
2435 => "00010000",
2436 => "00010000",
2437 => "00010000",
2438 => "00010000",
2439 => "00010000",
2440 => "00010000",
2441 => "00010000",
2442 => "00010000",
2443 => "00010000",
2444 => "00010000",
2445 => "00010000",
2446 => "00010000",
2447 => "00010000",
2448 => "00010000",
2449 => "00010000",
2450 => "00010000",
2451 => "00010000",
2452 => "00001100",
2453 => "00010000",
2454 => "00001100",
2455 => "00010000",
2456 => "01010101",
2457 => "10111111",
2458 => "00000101",
2459 => "00000001",
2460 => "00000001",
2461 => "00000001",
2462 => "00100101",
2463 => "10010110",
2464 => "11011111",
2465 => "11011111",
2466 => "11011111",
2467 => "11011111",
2468 => "11011111",
2469 => "11011111",
2470 => "11011111",
2471 => "11011111",
2472 => "11011111",
2473 => "11011111",
2474 => "11011111",
2475 => "11011111",
2476 => "11011111",
2477 => "11011111",
2478 => "11011111",
2479 => "11011111",
2480 => "11011111",
2481 => "11011111",
2482 => "11011111",
2483 => "11011111",
2484 => "11011111",
2485 => "11011111",
2486 => "11011111",
2487 => "11011111",
2488 => "11011111",
2489 => "11011111",
2490 => "11011111",
2491 => "11011111",
2492 => "11011111",
2493 => "11011111",
2494 => "11011111",
2495 => "11011111",
2496 => "11011111",
2497 => "11011111",
2498 => "11011111",
2499 => "11011111",
2500 => "11011111",
2501 => "11011111",
2502 => "11011111",
2503 => "11011111",
2504 => "11011111",
2505 => "11011111",
2506 => "11011111",
2507 => "11011111",
2508 => "11011111",
2509 => "11011111",
2510 => "11011111",
2511 => "11011111",
2512 => "11011111",
2513 => "11011111",
2514 => "11011111",
2515 => "11011111",
2516 => "11011111",
2517 => "11011111",
2518 => "11011111",
2519 => "11011111",
2520 => "11011111",
2521 => "11011111",
2522 => "11011111",
2523 => "11011111",
2524 => "11011111",
2525 => "11011111",
2526 => "11011111",
2527 => "11011111",
2528 => "11011111",
2529 => "11011111",
2530 => "11011111",
2531 => "11011111",
2532 => "11011111",
2533 => "11011111",
2534 => "11011111",
2535 => "11011111",
2536 => "11011111",
2537 => "11011111",
2538 => "10010110",
2539 => "00000101",
2540 => "00000000",
2541 => "00000001",
2542 => "00000001",
2543 => "00000001",
2544 => "00000000",
2545 => "00000000",
2546 => "00000000",
2547 => "00000000",
2548 => "00000000",
2549 => "00000000",
2550 => "00000000",
2551 => "00000000",
2552 => "00000000",
2553 => "00000000",
2554 => "00000000",
2555 => "00000000",
2556 => "00000000",
2557 => "00000000",
2558 => "00000000",
2559 => "00000000",
2560 => "00000000",
2561 => "00000000",
2562 => "00000000",
2563 => "00000000",
2564 => "00000000",
2565 => "00000000",
2566 => "00000000",
2567 => "00000000",
2568 => "00000000",
2569 => "00000000",
2570 => "00000000",
2571 => "00000000",
2572 => "00000000",
2573 => "00000000",
2574 => "00000000",
2575 => "00000000",
2576 => "00000000",
2577 => "00000000",
2578 => "00000000",
2579 => "00000000",
2580 => "00000000",
2581 => "00000000",
2582 => "00000000",
2583 => "00000000",
2584 => "00000000",
2585 => "00000000",
2586 => "00000000",
2587 => "00000000",
2588 => "00000000",
2589 => "00000000",
2590 => "00000000",
2591 => "00000000",
2592 => "00000000",
2593 => "00000000",
2594 => "00000000",
2595 => "00000000",
2596 => "00000000",
2597 => "00000000",
2598 => "00000000",
2599 => "00000000",
2600 => "00000000",
2601 => "00000000",
2602 => "00000000",
2603 => "00000000",
2604 => "00000000",
2605 => "00000000",
2606 => "00000000",
2607 => "00000000",
2608 => "00000000",
2609 => "00000000",
2610 => "00000000",
2611 => "00000000",
2612 => "00000000",
2613 => "00000000",
2614 => "00000000",
2615 => "00000000",
2616 => "00000000",
2617 => "00000000",
2618 => "00000000",
2619 => "00000000",
2620 => "00000001",
2621 => "00000001",
2622 => "00000001",
2623 => "00000001");
begin

    process(clk)
    begin
    
        if rising_edge(clk) then
                dout <= green(to_integer(unsigned(addr)));
        end if;
    end process;

end Behavioral;


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity SeverityAxis is
    port(clk, rst: in std_logic;
         addr: in std_logic_vector(10 downto 0);
         dout: out std_logic_vector(7 downto 0));
end SeverityAxis;

architecture Behavioral of SeverityAxis is

    type mem is array (0 to 1169) of std_logic_vector(7 downto 0);
    signal Class: mem := (
        0 => "00000000",
        1 => "00000000",
        2 => "00000000",
        3 => "00000000",
        4 => "00000000",
        5 => "00000000",
        6 => "00000000",
        7 => "00000000",
        8 => "00100100",
        9 => "11011010",
        10 => "01001000",
        11 => "00000000",
        12 => "00000000",
        13 => "00000000",
        14 => "00000000",
        15 => "00000000",
        16 => "00000000",
        17 => "00000000",
        18 => "00000000",
        19 => "00000000",
        20 => "00000000",
        21 => "00100100",
        22 => "11011010",
        23 => "01001000",
        24 => "00000000",
        25 => "00000000",
        26 => "00000000",
        27 => "10010001",
        28 => "11111111",
        29 => "11111111",
        30 => "11111111",
        31 => "11111111",
        32 => "11111111",
        33 => "11111111",
        34 => "11111111",
        35 => "11111111",
        36 => "01001000",
        37 => "00000000",
        38 => "00000000",
        39 => "00000000",
        40 => "10010001",
        41 => "10110110",
        42 => "00000000",
        43 => "00000000",
        44 => "00000000",
        45 => "00000000",
        46 => "00000000",
        47 => "00100100",
        48 => "11011010",
        49 => "01001000",
        50 => "00000000",
        51 => "00000000",
        52 => "00000000",
        53 => "10010001",
        54 => "10110110",
        55 => "00000000",
        56 => "00000000",
        57 => "00000000",
        58 => "00000000",
        59 => "00000000",
        60 => "00100100",
        61 => "11011010",
        62 => "01001000",
        63 => "00000000",
        64 => "00000000",
        65 => "00000000",
        66 => "00000000",
        67 => "00000000",
        68 => "00000000",
        69 => "00000000",
        70 => "00000000",
        71 => "00000000",
        72 => "00000000",
        73 => "00000000",
        74 => "00000000",
        75 => "00000000",
        76 => "00000000",
        77 => "00000000",
        78 => "00000000",
        79 => "00000000",
        80 => "00000000",
        81 => "00000000",
        82 => "01101101",
        83 => "11111111",
        84 => "11111111",
        85 => "10010001",
        86 => "01001000",
        87 => "11011010",
        88 => "00100100",
        89 => "00000000",
        90 => "00000000",
        91 => "00000000",
        92 => "00000000",
        93 => "00000000",
        94 => "00100100",
        95 => "11011010",
        96 => "01101101",
        97 => "10110110",
        98 => "10010001",
        99 => "00100100",
        100 => "11011010",
        101 => "01001000",
        102 => "00000000",
        103 => "00000000",
        104 => "00000000",
        105 => "00000000",
        106 => "00000000",
        107 => "01001000",
        108 => "11011010",
        109 => "00100100",
        110 => "10110110",
        111 => "10010001",
        112 => "00100100",
        113 => "11011010",
        114 => "01001000",
        115 => "00000000",
        116 => "00000000",
        117 => "00000000",
        118 => "00000000",
        119 => "00000000",
        120 => "00100100",
        121 => "11011011",
        122 => "10010001",
        123 => "10110110",
        124 => "10010001",
        125 => "10010001",
        126 => "11011011",
        127 => "00100100",
        128 => "00000000",
        129 => "00000000",
        130 => "00000000",
        131 => "00000000",
        132 => "00000000",
        133 => "00000000",
        134 => "00100100",
        135 => "11011011",
        136 => "11111111",
        137 => "11111111",
        138 => "11111111",
        139 => "01001000",
        140 => "00000000",
        141 => "00000000",
        142 => "00000000",
        143 => "00000000",
        144 => "00000000",
        145 => "00000000",
        146 => "00000000",
        147 => "00000000",
        148 => "00000000",
        149 => "00000000",
        150 => "00000000",
        151 => "00000000",
        152 => "00000000",
        153 => "00000000",
        154 => "00000000",
        155 => "00000000",
        156 => "00000000",
        157 => "00000000",
        158 => "00000000",
        159 => "00000000",
        160 => "00000000",
        161 => "00000000",
        162 => "00000000",
        163 => "00000000",
        164 => "00000000",
        165 => "00000000",
        166 => "00000000",
        167 => "00000000",
        168 => "00000000",
        169 => "00000000",
        170 => "00000000",
        171 => "00000000",
        172 => "00100100",
        173 => "11011011",
        174 => "11111111",
        175 => "11011010",
        176 => "00000000",
        177 => "00000000",
        178 => "00000000",
        179 => "00000000",
        180 => "00000000",
        181 => "00000000",
        182 => "00000000",
        183 => "00000000",
        184 => "00000000",
        185 => "00000000",
        186 => "00000000",
        187 => "00000000",
        188 => "10010001",
        189 => "11111111",
        190 => "11111111",
        191 => "10010001",
        192 => "00000000",
        193 => "00000000",
        194 => "00000000",
        195 => "00000000",
        196 => "00000000",
        197 => "00000000",
        198 => "00000000",
        199 => "00000000",
        200 => "00000000",
        201 => "00000000",
        202 => "00000000",
        203 => "00000000",
        204 => "10110110",
        205 => "01001000",
        206 => "00000000",
        207 => "00000000",
        208 => "00000000",
        209 => "00000000",
        210 => "00000000",
        211 => "00000000",
        212 => "00000000",
        213 => "00000000",
        214 => "10010001",
        215 => "11111111",
        216 => "11111111",
        217 => "10010001",
        218 => "00000000",
        219 => "00000000",
        220 => "00000000",
        221 => "00000000",
        222 => "00000000",
        223 => "00000000",
        224 => "00100100",
        225 => "11011011",
        226 => "11111111",
        227 => "11011010",
        228 => "00000000",
        229 => "00000000",
        230 => "00000000",
        231 => "00000000",
        232 => "00000000",
        233 => "00000000",
        234 => "00000000",
        235 => "00000000",
        236 => "00000000",
        237 => "00000000",
        238 => "00000000",
        239 => "00000000",
        240 => "00000000",
        241 => "00000000",
        242 => "00000000",
        243 => "00000000",
        244 => "00000000",
        245 => "00000000",
        246 => "00000000",
        247 => "00000000",
        248 => "00000000",
        249 => "00000000",
        250 => "00000000",
        251 => "01101101",
        252 => "11111111",
        253 => "11111111",
        254 => "10010001",
        255 => "01001000",
        256 => "11011010",
        257 => "00100100",
        258 => "00000000",
        259 => "00000000",
        260 => "00000000",
        261 => "00000000",
        262 => "00000000",
        263 => "00100100",
        264 => "11011010",
        265 => "01101101",
        266 => "10110110",
        267 => "10010001",
        268 => "00100100",
        269 => "11011010",
        270 => "01001000",
        271 => "00000000",
        272 => "00000000",
        273 => "00000000",
        274 => "00000000",
        275 => "00000000",
        276 => "01001000",
        277 => "11011010",
        278 => "00100100",
        279 => "10110110",
        280 => "10010001",
        281 => "00100100",
        282 => "11011010",
        283 => "01001000",
        284 => "00000000",
        285 => "00000000",
        286 => "00000000",
        287 => "00000000",
        288 => "00000000",
        289 => "00100100",
        290 => "11011011",
        291 => "10010001",
        292 => "10110110",
        293 => "10010001",
        294 => "10010001",
        295 => "11011011",
        296 => "00100100",
        297 => "00000000",
        298 => "00000000",
        299 => "00000000",
        300 => "00000000",
        301 => "00000000",
        302 => "00000000",
        303 => "00100100",
        304 => "11011011",
        305 => "11111111",
        306 => "11111111",
        307 => "11111111",
        308 => "01001000",
        309 => "00000000",
        310 => "00000000",
        311 => "00000000",
        312 => "00000000",
        313 => "00000000",
        314 => "00000000",
        315 => "00000000",
        316 => "00000000",
        317 => "00000000",
        318 => "00000000",
        319 => "00000000",
        320 => "00000000",
        321 => "00000000",
        322 => "00000000",
        323 => "00000000",
        324 => "00000000",
        325 => "00000000",
        326 => "00000000",
        327 => "00000000",
        328 => "00000000",
        329 => "00000000",
        330 => "00000000",
        331 => "00000000",
        332 => "00000000",
        333 => "00000000",
        334 => "00000000",
        335 => "00000000",
        336 => "00000000",
        337 => "00000000",
        338 => "00000000",
        339 => "00000000",
        340 => "00000000",
        341 => "00000000",
        342 => "00000000",
        343 => "00000000",
        344 => "00000000",
        345 => "00000000",
        346 => "00000000",
        347 => "00000000",
        348 => "00000000",
        349 => "00000000",
        350 => "00000000",
        351 => "00000000",
        352 => "00000000",
        353 => "00000000",
        354 => "00000000",
        355 => "00000000",
        356 => "00000000",
        357 => "00000000",
        358 => "00000000",
        359 => "00100100",
        360 => "11011010",
        361 => "01001000",
        362 => "00000000",
        363 => "00000000",
        364 => "00000000",
        365 => "00000000",
        366 => "00000000",
        367 => "00000000",
        368 => "00000000",
        369 => "00000000",
        370 => "00000000",
        371 => "00000000",
        372 => "00100100",
        373 => "11011010",
        374 => "01001000",
        375 => "00000000",
        376 => "00000000",
        377 => "00000000",
        378 => "00000000",
        379 => "00000000",
        380 => "00000000",
        381 => "00000000",
        382 => "00000000",
        383 => "00000000",
        384 => "00000000",
        385 => "00100100",
        386 => "11011010",
        387 => "01001000",
        388 => "00000000",
        389 => "00000000",
        390 => "00000000",
        391 => "00000000",
        392 => "11011010",
        393 => "11111111",
        394 => "11111111",
        395 => "11111111",
        396 => "11111111",
        397 => "11111111",
        398 => "11111111",
        399 => "11111111",
        400 => "01001000",
        401 => "00000000",
        402 => "00000000",
        403 => "00000000",
        404 => "00000000",
        405 => "00000000",
        406 => "00000000",
        407 => "00000000",
        408 => "00000000",
        409 => "00000000",
        410 => "00000000",
        411 => "00000000",
        412 => "00000000",
        413 => "00000000",
        414 => "00000000",
        415 => "00000000",
        416 => "00000000",
        417 => "00000000",
        418 => "00000000",
        419 => "00000000",
        420 => "00000000",
        421 => "00000000",
        422 => "00000000",
        423 => "00000000",
        424 => "00000000",
        425 => "00000000",
        426 => "00000000",
        427 => "00000000",
        428 => "00000000",
        429 => "00000000",
        430 => "00000000",
        431 => "00000000",
        432 => "00000000",
        433 => "00000000",
        434 => "00000000",
        435 => "00000000",
        436 => "00000000",
        437 => "00000000",
        438 => "00000000",
        439 => "00000000",
        440 => "00000000",
        441 => "00000000",
        442 => "00000000",
        443 => "00000000",
        444 => "00000000",
        445 => "00000000",
        446 => "00000000",
        447 => "00000000",
        448 => "00000000",
        449 => "00000000",
        450 => "00000000",
        451 => "00000000",
        452 => "00000000",
        453 => "00000000",
        454 => "00000000",
        455 => "00000000",
        456 => "00000000",
        457 => "00000000",
        458 => "00000000",
        459 => "00000000",
        460 => "00000000",
        461 => "00000000",
        462 => "00000000",
        463 => "00000000",
        464 => "00000000",
        465 => "00000000",
        466 => "00000000",
        467 => "00000000",
        468 => "00000000",
        469 => "00000000",
        470 => "00000000",
        471 => "00000000",
        472 => "00000000",
        473 => "00000000",
        474 => "00000000",
        475 => "00000000",
        476 => "00000000",
        477 => "00000000",
        478 => "00000000",
        479 => "00000000",
        480 => "00000000",
        481 => "00000000",
        482 => "00000000",
        483 => "00000000",
        484 => "00000000",
        485 => "00000000",
        486 => "00000000",
        487 => "00000000",
        488 => "00000000",
        489 => "00000000",
        490 => "00000000",
        491 => "00000000",
        492 => "00000000",
        493 => "00000000",
        494 => "00000000",
        495 => "00000000",
        496 => "00000000",
        497 => "00000000",
        498 => "00000000",
        499 => "00000000",
        500 => "00000000",
        501 => "00000000",
        502 => "00000000",
        503 => "00000000",
        504 => "00000000",
        505 => "00000000",
        506 => "00000000",
        507 => "00000000",
        508 => "00000000",
        509 => "00000000",
        510 => "00100100",
        511 => "11011011",
        512 => "11111111",
        513 => "01101101",
        514 => "00000000",
        515 => "00000000",
        516 => "00000000",
        517 => "00000000",
        518 => "00000000",
        519 => "00000000",
        520 => "00000000",
        521 => "00000000",
        522 => "00000000",
        523 => "00000000",
        524 => "00000000",
        525 => "00100100",
        526 => "11011011",
        527 => "11111111",
        528 => "10110110",
        529 => "00000000",
        530 => "00000000",
        531 => "00000000",
        532 => "00000000",
        533 => "00000000",
        534 => "00000000",
        535 => "00000000",
        536 => "00000000",
        537 => "00000000",
        538 => "00000000",
        539 => "00000000",
        540 => "00000000",
        541 => "10110110",
        542 => "11111111",
        543 => "10110110",
        544 => "00000000",
        545 => "00000000",
        546 => "00000000",
        547 => "00000000",
        548 => "00000000",
        549 => "00000000",
        550 => "00000000",
        551 => "00000000",
        552 => "10110110",
        553 => "11111111",
        554 => "11111111",
        555 => "01001000",
        556 => "10110110",
        557 => "11011010",
        558 => "00000000",
        559 => "00000000",
        560 => "00000000",
        561 => "00000000",
        562 => "00100100",
        563 => "11011011",
        564 => "11111111",
        565 => "10110110",
        566 => "00000000",
        567 => "00000000",
        568 => "00000000",
        569 => "00100100",
        570 => "11011010",
        571 => "01001000",
        572 => "00000000",
        573 => "00000000",
        574 => "00000000",
        575 => "00000000",
        576 => "00000000",
        577 => "00000000",
        578 => "00000000",
        579 => "00000000",
        580 => "00000000",
        581 => "00000000",
        582 => "01001000",
        583 => "11011011",
        584 => "01001000",
        585 => "00000000",
        586 => "00000000",
        587 => "00000000",
        588 => "00000000",
        589 => "00000000",
        590 => "00000000",
        591 => "00000000",
        592 => "00000000",
        593 => "00000000",
        594 => "00000000",
        595 => "00000000",
        596 => "00000000",
        597 => "00000000",
        598 => "00000000",
        599 => "00000000",
        600 => "00000000",
        601 => "00000000",
        602 => "00000000",
        603 => "00000000",
        604 => "00000000",
        605 => "00000000",
        606 => "00000000",
        607 => "00000000",
        608 => "00000000",
        609 => "00000000",
        610 => "00000000",
        611 => "00000000",
        612 => "00000000",
        613 => "00000000",
        614 => "00100100",
        615 => "11011010",
        616 => "01001000",
        617 => "00000000",
        618 => "00000000",
        619 => "01001000",
        620 => "11011011",
        621 => "01001000",
        622 => "00000000",
        623 => "00000000",
        624 => "00000000",
        625 => "00000000",
        626 => "00000000",
        627 => "00100100",
        628 => "11011010",
        629 => "01001000",
        630 => "00000000",
        631 => "00000000",
        632 => "00100100",
        633 => "11011010",
        634 => "01001000",
        635 => "00000000",
        636 => "00000000",
        637 => "00000000",
        638 => "00000000",
        639 => "11011010",
        640 => "11111111",
        641 => "11111111",
        642 => "11111111",
        643 => "11111111",
        644 => "11111111",
        645 => "11111111",
        646 => "11011011",
        647 => "00100100",
        648 => "00000000",
        649 => "00000000",
        650 => "00000000",
        651 => "00000000",
        652 => "00000000",
        653 => "00100100",
        654 => "11011010",
        655 => "01001000",
        656 => "00000000",
        657 => "00000000",
        658 => "00000000",
        659 => "00000000",
        660 => "00000000",
        661 => "00000000",
        662 => "00000000",
        663 => "00000000",
        664 => "00000000",
        665 => "00000000",
        666 => "00100100",
        667 => "11011010",
        668 => "01001000",
        669 => "00000000",
        670 => "00000000",
        671 => "00000000",
        672 => "00000000",
        673 => "00000000",
        674 => "00000000",
        675 => "00000000",
        676 => "00000000",
        677 => "00000000",
        678 => "00000000",
        679 => "00000000",
        680 => "00000000",
        681 => "00000000",
        682 => "00000000",
        683 => "00000000",
        684 => "00100100",
        685 => "11011010",
        686 => "01001000",
        687 => "00000000",
        688 => "00000000",
        689 => "00000000",
        690 => "01001000",
        691 => "11011011",
        692 => "01001000",
        693 => "00000000",
        694 => "00000000",
        695 => "00000000",
        696 => "00000000",
        697 => "00100100",
        698 => "11011010",
        699 => "01001000",
        700 => "00000000",
        701 => "00000000",
        702 => "00000000",
        703 => "01101101",
        704 => "11111111",
        705 => "10010001",
        706 => "11011011",
        707 => "11111111",
        708 => "11111111",
        709 => "11111111",
        710 => "11111111",
        711 => "11111111",
        712 => "01001000",
        713 => "00000000",
        714 => "00000000",
        715 => "00000000",
        716 => "00000000",
        717 => "00000000",
        718 => "00100100",
        719 => "11011010",
        720 => "01001000",
        721 => "00000000",
        722 => "00000000",
        723 => "00100100",
        724 => "11011010",
        725 => "01001000",
        726 => "00000000",
        727 => "00000000",
        728 => "00000000",
        729 => "00000000",
        730 => "00000000",
        731 => "00100100",
        732 => "11011010",
        733 => "01001000",
        734 => "00000000",
        735 => "00000000",
        736 => "00100100",
        737 => "11011010",
        738 => "01001000",
        739 => "00000000",
        740 => "00000000",
        741 => "00000000",
        742 => "00000000",
        743 => "00000000",
        744 => "00000000",
        745 => "00000000",
        746 => "00000000",
        747 => "00000000",
        748 => "00000000",
        749 => "00000000",
        750 => "00000000",
        751 => "00000000",
        752 => "00000000",
        753 => "00000000",
        754 => "00000000",
        755 => "00000000",
        756 => "00000000",
        757 => "00000000",
        758 => "00000000",
        759 => "00000000",
        760 => "00000000",
        761 => "00000000",
        762 => "00000000",
        763 => "00000000",
        764 => "00000000",
        765 => "00000000",
        766 => "00000000",
        767 => "00000000",
        768 => "00000000",
        769 => "00000000",
        770 => "00000000",
        771 => "10110110",
        772 => "11111111",
        773 => "10010001",
        774 => "00000000",
        775 => "00000000",
        776 => "00000000",
        777 => "00000000",
        778 => "00000000",
        779 => "00000000",
        780 => "00000000",
        781 => "00000000",
        782 => "00000000",
        783 => "01001000",
        784 => "11011011",
        785 => "01001000",
        786 => "00000000",
        787 => "00000000",
        788 => "00000000",
        789 => "00000000",
        790 => "00000000",
        791 => "00000000",
        792 => "00000000",
        793 => "00000000",
        794 => "00000000",
        795 => "00000000",
        796 => "00100100",
        797 => "11011010",
        798 => "01001000",
        799 => "00000000",
        800 => "00000000",
        801 => "00000000",
        802 => "00000000",
        803 => "00000000",
        804 => "00000000",
        805 => "00000000",
        806 => "00000000",
        807 => "00000000",
        808 => "00000000",
        809 => "00000000",
        810 => "10010001",
        811 => "11011010",
        812 => "00000000",
        813 => "00000000",
        814 => "00000000",
        815 => "00000000",
        816 => "00000000",
        817 => "00000000",
        818 => "00000000",
        819 => "00000000",
        820 => "00000000",
        821 => "00000000",
        822 => "00100100",
        823 => "11011011",
        824 => "11111111",
        825 => "11111111",
        826 => "11111111",
        827 => "11111111",
        828 => "11111111",
        829 => "01001000",
        830 => "00000000",
        831 => "00000000",
        832 => "00000000",
        833 => "00000000",
        834 => "00000000",
        835 => "00000000",
        836 => "00000000",
        837 => "00000000",
        838 => "00000000",
        839 => "00000000",
        840 => "00000000",
        841 => "00000000",
        842 => "00000000",
        843 => "00000000",
        844 => "00000000",
        845 => "00000000",
        846 => "00000000",
        847 => "00000000",
        848 => "00000000",
        849 => "00000000",
        850 => "00000000",
        851 => "00000000",
        852 => "00000000",
        853 => "00000000",
        854 => "00000000",
        855 => "00000000",
        856 => "00000000",
        857 => "00000000",
        858 => "00000000",
        859 => "00000000",
        860 => "00000000",
        861 => "00000000",
        862 => "01101101",
        863 => "11111111",
        864 => "11111111",
        865 => "10010001",
        866 => "01001000",
        867 => "11011010",
        868 => "00100100",
        869 => "00000000",
        870 => "00000000",
        871 => "00000000",
        872 => "00000000",
        873 => "00000000",
        874 => "00100100",
        875 => "11011010",
        876 => "01101101",
        877 => "10110110",
        878 => "10010001",
        879 => "00100100",
        880 => "11011010",
        881 => "01001000",
        882 => "00000000",
        883 => "00000000",
        884 => "00000000",
        885 => "00000000",
        886 => "00000000",
        887 => "01001000",
        888 => "11011010",
        889 => "00100100",
        890 => "10110110",
        891 => "10010001",
        892 => "00100100",
        893 => "11011010",
        894 => "01001000",
        895 => "00000000",
        896 => "00000000",
        897 => "00000000",
        898 => "00000000",
        899 => "00000000",
        900 => "00100100",
        901 => "11011011",
        902 => "10010001",
        903 => "10110110",
        904 => "10010001",
        905 => "10010001",
        906 => "11011011",
        907 => "00100100",
        908 => "00000000",
        909 => "00000000",
        910 => "00000000",
        911 => "00000000",
        912 => "00000000",
        913 => "00000000",
        914 => "00100100",
        915 => "11011011",
        916 => "11111111",
        917 => "11111111",
        918 => "11111111",
        919 => "01001000",
        920 => "00000000",
        921 => "00000000",
        922 => "00000000",
        923 => "00000000",
        924 => "00000000",
        925 => "00000000",
        926 => "00000000",
        927 => "00000000",
        928 => "00000000",
        929 => "00000000",
        930 => "00000000",
        931 => "00000000",
        932 => "00000000",
        933 => "00000000",
        934 => "00000000",
        935 => "00000000",
        936 => "00000000",
        937 => "00000000",
        938 => "00000000",
        939 => "00100100",
        940 => "11011011",
        941 => "11111111",
        942 => "11011010",
        943 => "00000000",
        944 => "00000000",
        945 => "00000000",
        946 => "00000000",
        947 => "00000000",
        948 => "00000000",
        949 => "00000000",
        950 => "00000000",
        951 => "00000000",
        952 => "00000000",
        953 => "00000000",
        954 => "00000000",
        955 => "10010001",
        956 => "11111111",
        957 => "11111111",
        958 => "10010001",
        959 => "00000000",
        960 => "00000000",
        961 => "00000000",
        962 => "00000000",
        963 => "00000000",
        964 => "00000000",
        965 => "00000000",
        966 => "00000000",
        967 => "00000000",
        968 => "00000000",
        969 => "00000000",
        970 => "00000000",
        971 => "10110110",
        972 => "01001000",
        973 => "00000000",
        974 => "00000000",
        975 => "00000000",
        976 => "00000000",
        977 => "00000000",
        978 => "00000000",
        979 => "00000000",
        980 => "00000000",
        981 => "10010001",
        982 => "11111111",
        983 => "11111111",
        984 => "10010001",
        985 => "00000000",
        986 => "00000000",
        987 => "00000000",
        988 => "00000000",
        989 => "00000000",
        990 => "00000000",
        991 => "00100100",
        992 => "11011011",
        993 => "11111111",
        994 => "11011010",
        995 => "00000000",
        996 => "00000000",
        997 => "00000000",
        998 => "00000000",
        999 => "00000000",
        1000 => "00000000",
        1001 => "00000000",
        1002 => "00000000",
        1003 => "00000000",
        1004 => "00000000",
        1005 => "00000000",
        1006 => "00000000",
        1007 => "00000000",
        1008 => "00000000",
        1009 => "00000000",
        1010 => "00000000",
        1011 => "00000000",
        1012 => "00000000",
        1013 => "00000000",
        1014 => "00000000",
        1015 => "00000000",
        1016 => "00000000",
        1017 => "00000000",
        1018 => "00000000",
        1019 => "00000000",
        1020 => "00000000",
        1021 => "00000000",
        1022 => "00000000",
        1023 => "00000000",
        1024 => "00000000",
        1025 => "00000000",
        1026 => "00000000",
        1027 => "00000000",
        1028 => "00000000",
        1029 => "00000000",
        1030 => "00000000",
        1031 => "01101101",
        1032 => "11111111",
        1033 => "11111111",
        1034 => "10010001",
        1035 => "01001000",
        1036 => "11011010",
        1037 => "00100100",
        1038 => "00000000",
        1039 => "00000000",
        1040 => "00000000",
        1041 => "00000000",
        1042 => "00000000",
        1043 => "00100100",
        1044 => "11011010",
        1045 => "01101101",
        1046 => "10110110",
        1047 => "10010001",
        1048 => "00100100",
        1049 => "11011010",
        1050 => "01001000",
        1051 => "00000000",
        1052 => "00000000",
        1053 => "00000000",
        1054 => "00000000",
        1055 => "00000000",
        1056 => "01001000",
        1057 => "11011010",
        1058 => "00100100",
        1059 => "10110110",
        1060 => "10010001",
        1061 => "00100100",
        1062 => "11011010",
        1063 => "01001000",
        1064 => "00000000",
        1065 => "00000000",
        1066 => "00000000",
        1067 => "00000000",
        1068 => "00000000",
        1069 => "00100100",
        1070 => "11011011",
        1071 => "10010001",
        1072 => "10110110",
        1073 => "10010001",
        1074 => "10010001",
        1075 => "11011011",
        1076 => "00100100",
        1077 => "00000000",
        1078 => "00000000",
        1079 => "00000000",
        1080 => "00000000",
        1081 => "00000000",
        1082 => "00000000",
        1083 => "00100100",
        1084 => "11011011",
        1085 => "11111111",
        1086 => "11111111",
        1087 => "11111111",
        1088 => "01001000",
        1089 => "00000000",
        1090 => "00000000",
        1091 => "00000000",
        1092 => "00000000",
        1093 => "00000000",
        1094 => "00000000",
        1095 => "00000000",
        1096 => "00000000",
        1097 => "00000000",
        1098 => "00000000",
        1099 => "00000000",
        1100 => "00000000",
        1101 => "00000000",
        1102 => "00000000",
        1103 => "00000000",
        1104 => "00000000",
        1105 => "00000000",
        1106 => "01001000",
        1107 => "11011011",
        1108 => "01001000",
        1109 => "00000000",
        1110 => "00000000",
        1111 => "11011010",
        1112 => "11111111",
        1113 => "11111111",
        1114 => "10010001",
        1115 => "00000000",
        1116 => "00000000",
        1117 => "00000000",
        1118 => "00000000",
        1119 => "01001000",
        1120 => "11011010",
        1121 => "00100100",
        1122 => "00000000",
        1123 => "01101101",
        1124 => "11011011",
        1125 => "01001000",
        1126 => "01101101",
        1127 => "11011010",
        1128 => "00100100",
        1129 => "00000000",
        1130 => "00000000",
        1131 => "00000000",
        1132 => "01001000",
        1133 => "11011010",
        1134 => "00100100",
        1135 => "00000000",
        1136 => "11011010",
        1137 => "10110110",
        1138 => "00000000",
        1139 => "00100100",
        1140 => "11011010",
        1141 => "01001000",
        1142 => "00000000",
        1143 => "00000000",
        1144 => "00000000",
        1145 => "00000000",
        1146 => "11011010",
        1147 => "10010001",
        1148 => "01101101",
        1149 => "11011011",
        1150 => "01001000",
        1151 => "00000000",
        1152 => "00100100",
        1153 => "11011010",
        1154 => "01001000",
        1155 => "00000000",
        1156 => "00000000",
        1157 => "00000000",
        1158 => "00000000",
        1159 => "01101101",
        1160 => "11111111",
        1161 => "11111111",
        1162 => "10010001",
        1163 => "00000000",
        1164 => "00000000",
        1165 => "01101101",
        1166 => "11011010",
        1167 => "00100100",
        1168 => "00000000",
        1169 => "00000000");

begin

    process(clk)
    begin
    
        if rising_edge(clk) then
            if rst = '1' then
                Class <= (others => (others => '0'));
            else
                dout <= Class(to_integer(unsigned(addr)));
            end if;
        end if;
    end process;

end Behavioral;

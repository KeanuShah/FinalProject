
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity FreqAxis is
     port(clk, rst: in std_logic;
         addr: in std_logic_vector(10 downto 0);
         dout: out std_logic_vector(7 downto 0));
end FreqAxis;

architecture Behavioral of FreqAxis is

    type mem is array (0 to 1067) of std_logic_vector(7 downto 0);
    signal Freq: mem := (
        0 => "00000000",
        1 => "00000000",
        2 => "01001000",
        3 => "11111111",
        4 => "11111111",
        5 => "11111111",
        6 => "11111111",
        7 => "11111111",
        8 => "01101101",
        9 => "00000000",
        10 => "00000000",
        11 => "00000000",
        12 => "00000000",
        13 => "11011010",
        14 => "11111111",
        15 => "01101101",
        16 => "00000000",
        17 => "00000000",
        18 => "00000000",
        19 => "00100100",
        20 => "11011011",
        21 => "11111111",
        22 => "01001000",
        23 => "00000000",
        24 => "11011010",
        25 => "10110110",
        26 => "00000000",
        27 => "00000000",
        28 => "00000000",
        29 => "00000000",
        30 => "00000000",
        31 => "00000000",
        32 => "00000000",
        33 => "01101101",
        34 => "11011011",
        35 => "01001000",
        36 => "00000000",
        37 => "00000000",
        38 => "00000000",
        39 => "00000000",
        40 => "00000000",
        41 => "00000000",
        42 => "00000000",
        43 => "00000000",
        44 => "00000000",
        45 => "00000000",
        46 => "00000000",
        47 => "00000000",
        48 => "00000000",
        49 => "00000000",
        50 => "00000000",
        51 => "00000000",
        52 => "00000000",
        53 => "00000000",
        54 => "00000000",
        55 => "00000000",
        56 => "00000000",
        57 => "00000000",
        58 => "00000000",
        59 => "00000000",
        60 => "00000000",
        61 => "00000000",
        62 => "00100100",
        63 => "11011010",
        64 => "01101101",
        65 => "00000000",
        66 => "00000000",
        67 => "00100100",
        68 => "11011010",
        69 => "01001000",
        70 => "00000000",
        71 => "00000000",
        72 => "00000000",
        73 => "00000000",
        74 => "00100100",
        75 => "11011010",
        76 => "11111111",
        77 => "10110110",
        78 => "00000000",
        79 => "00100100",
        80 => "11011010",
        81 => "01001000",
        82 => "00000000",
        83 => "00000000",
        84 => "00000000",
        85 => "00000000",
        86 => "00100100",
        87 => "11011010",
        88 => "01001000",
        89 => "10110110",
        90 => "11011010",
        91 => "00100100",
        92 => "11011010",
        93 => "01001000",
        94 => "00000000",
        95 => "00000000",
        96 => "00000000",
        97 => "00000000",
        98 => "00100100",
        99 => "11011010",
        100 => "01001000",
        101 => "00000000",
        102 => "10010001",
        103 => "11111111",
        104 => "11011011",
        105 => "01001000",
        106 => "00000000",
        107 => "00000000",
        108 => "00000000",
        109 => "00000000",
        110 => "00100100",
        111 => "11011010",
        112 => "01001000",
        113 => "00000000",
        114 => "00000000",
        115 => "01001000",
        116 => "11011011",
        117 => "01001000",
        118 => "00000000",
        119 => "00000000",
        120 => "00000000",
        121 => "00000000",
        122 => "00000000",
        123 => "00000000",
        124 => "00000000",
        125 => "00000000",
        126 => "00000000",
        127 => "00000000",
        128 => "00000000",
        129 => "00000000",
        130 => "00000000",
        131 => "00000000",
        132 => "00000000",
        133 => "00000000",
        134 => "00000000",
        135 => "00000000",
        136 => "00000000",
        137 => "00000000",
        138 => "00000000",
        139 => "00000000",
        140 => "00000000",
        141 => "00000000",
        142 => "00000000",
        143 => "00000000",
        144 => "00000000",
        145 => "11011010",
        146 => "11111111",
        147 => "11111111",
        148 => "11111111",
        149 => "11111111",
        150 => "11111111",
        151 => "11111111",
        152 => "11111111",
        153 => "01001000",
        154 => "00000000",
        155 => "00000000",
        156 => "00000000",
        157 => "00000000",
        158 => "00000000",
        159 => "00000000",
        160 => "10110110",
        161 => "10110110",
        162 => "00000000",
        163 => "00000000",
        164 => "00000000",
        165 => "00000000",
        166 => "00000000",
        167 => "00000000",
        168 => "00000000",
        169 => "00000000",
        170 => "00000000",
        171 => "00000000",
        172 => "10110110",
        173 => "10110110",
        174 => "00000000",
        175 => "00000000",
        176 => "00000000",
        177 => "00000000",
        178 => "00000000",
        179 => "00000000",
        180 => "00000000",
        181 => "00000000",
        182 => "00000000",
        183 => "00000000",
        184 => "10110110",
        185 => "10110110",
        186 => "00000000",
        187 => "00000000",
        188 => "00000000",
        189 => "00000000",
        190 => "00000000",
        191 => "00000000",
        192 => "00000000",
        193 => "11011010",
        194 => "11111111",
        195 => "11111111",
        196 => "11111111",
        197 => "11111111",
        198 => "11111111",
        199 => "11111111",
        200 => "11111111",
        201 => "01001000",
        202 => "00000000",
        203 => "00000000",
        204 => "00000000",
        205 => "00000000",
        206 => "00000000",
        207 => "00000000",
        208 => "00000000",
        209 => "00000000",
        210 => "00000000",
        211 => "00000000",
        212 => "00000000",
        213 => "00000000",
        214 => "00000000",
        215 => "00000000",
        216 => "00000000",
        217 => "00000000",
        218 => "00000000",
        219 => "00000000",
        220 => "00000000",
        221 => "00000000",
        222 => "00000000",
        223 => "00000000",
        224 => "00000000",
        225 => "00000000",
        226 => "00000000",
        227 => "00000000",
        228 => "11011010",
        229 => "10010001",
        230 => "00000000",
        231 => "00000000",
        232 => "00000000",
        233 => "00000000",
        234 => "00000000",
        235 => "00000000",
        236 => "00000000",
        237 => "01101101",
        238 => "11011011",
        239 => "01001000",
        240 => "00000000",
        241 => "11011010",
        242 => "11111111",
        243 => "01101101",
        244 => "00000000",
        245 => "00000000",
        246 => "00000000",
        247 => "00100100",
        248 => "11011011",
        249 => "11111111",
        250 => "01001000",
        251 => "00000000",
        252 => "00000000",
        253 => "00000000",
        254 => "01001000",
        255 => "11111111",
        256 => "11111111",
        257 => "11111111",
        258 => "11111111",
        259 => "11111111",
        260 => "10010001",
        261 => "00000000",
        262 => "00000000",
        263 => "00000000",
        264 => "00000000",
        265 => "00000000",
        266 => "00000000",
        267 => "00000000",
        268 => "00000000",
        269 => "00000000",
        270 => "00000000",
        271 => "00000000",
        272 => "00000000",
        273 => "00000000",
        274 => "00000000",
        275 => "00000000",
        276 => "00000000",
        277 => "00000000",
        278 => "00000000",
        279 => "00000000",
        280 => "00000000",
        281 => "00000000",
        282 => "00000000",
        283 => "00000000",
        284 => "00000000",
        285 => "00000000",
        286 => "00000000",
        287 => "00000000",
        288 => "00000000",
        289 => "00000000",
        290 => "00000000",
        291 => "00000000",
        292 => "00000000",
        293 => "00000000",
        294 => "00000000",
        295 => "00000000",
        296 => "00000000",
        297 => "00000000",
        298 => "00000000",
        299 => "00000000",
        300 => "00000000",
        301 => "00000000",
        302 => "00000000",
        303 => "00000000",
        304 => "00000000",
        305 => "00000000",
        306 => "00000000",
        307 => "00000000",
        308 => "00000000",
        309 => "00000000",
        310 => "00000000",
        311 => "00000000",
        312 => "00000000",
        313 => "00000000",
        314 => "00000000",
        315 => "00000000",
        316 => "00000000",
        317 => "00000000",
        318 => "00000000",
        319 => "00000000",
        320 => "00000000",
        321 => "00000000",
        322 => "00000000",
        323 => "00000000",
        324 => "00000000",
        325 => "00000000",
        326 => "00000000",
        327 => "00000000",
        328 => "00000000",
        329 => "00000000",
        330 => "00000000",
        331 => "00000000",
        332 => "00000000",
        333 => "00000000",
        334 => "00000000",
        335 => "00000000",
        336 => "00000000",
        337 => "00000000",
        338 => "00000000",
        339 => "00000000",
        340 => "00000000",
        341 => "00000000",
        342 => "00000000",
        343 => "00000000",
        344 => "00000000",
        345 => "00000000",
        346 => "00000000",
        347 => "00000000",
        348 => "00000000",
        349 => "00000000",
        350 => "00000000",
        351 => "00000000",
        352 => "00000000",
        353 => "00000000",
        354 => "00000000",
        355 => "00000000",
        356 => "00000000",
        357 => "00000000",
        358 => "00000000",
        359 => "00000000",
        360 => "00000000",
        361 => "00000000",
        362 => "00000000",
        363 => "00000000",
        364 => "00000000",
        365 => "00000000",
        366 => "00000000",
        367 => "00000000",
        368 => "00000000",
        369 => "00000000",
        370 => "00000000",
        371 => "00000000",
        372 => "00000000",
        373 => "00000000",
        374 => "00000000",
        375 => "00000000",
        376 => "00000000",
        377 => "00000000",
        378 => "00000000",
        379 => "00000000",
        380 => "00000000",
        381 => "00000000",
        382 => "00000000",
        383 => "00000000",
        384 => "00000000",
        385 => "00000000",
        386 => "00100100",
        387 => "11011011",
        388 => "11111111",
        389 => "01101101",
        390 => "00000000",
        391 => "00000000",
        392 => "00000000",
        393 => "00000000",
        394 => "00000000",
        395 => "00000000",
        396 => "00000000",
        397 => "00000000",
        398 => "00000000",
        399 => "00000000",
        400 => "00100100",
        401 => "11011011",
        402 => "11111111",
        403 => "10110110",
        404 => "00000000",
        405 => "00000000",
        406 => "00000000",
        407 => "00000000",
        408 => "00000000",
        409 => "00000000",
        410 => "00000000",
        411 => "00000000",
        412 => "00000000",
        413 => "00000000",
        414 => "00000000",
        415 => "10110110",
        416 => "11111111",
        417 => "10110110",
        418 => "00000000",
        419 => "00000000",
        420 => "00000000",
        421 => "00000000",
        422 => "00000000",
        423 => "00000000",
        424 => "00000000",
        425 => "10110110",
        426 => "11111111",
        427 => "11111111",
        428 => "01001000",
        429 => "10110110",
        430 => "11011010",
        431 => "00000000",
        432 => "00000000",
        433 => "00000000",
        434 => "00100100",
        435 => "11011011",
        436 => "11111111",
        437 => "10110110",
        438 => "00000000",
        439 => "00000000",
        440 => "00000000",
        441 => "00100100",
        442 => "11011010",
        443 => "01001000",
        444 => "00000000",
        445 => "00000000",
        446 => "00000000",
        447 => "00000000",
        448 => "00000000",
        449 => "00000000",
        450 => "00000000",
        451 => "00000000",
        452 => "00000000",
        453 => "01001000",
        454 => "11011011",
        455 => "01001000",
        456 => "00000000",
        457 => "00000000",
        458 => "00100100",
        459 => "11011010",
        460 => "01101101",
        461 => "00000000",
        462 => "00000000",
        463 => "01101101",
        464 => "11011010",
        465 => "00100100",
        466 => "00000000",
        467 => "00000000",
        468 => "00000000",
        469 => "00000000",
        470 => "01001000",
        471 => "11011010",
        472 => "00100100",
        473 => "00000000",
        474 => "00000000",
        475 => "00100100",
        476 => "11011010",
        477 => "01001000",
        478 => "00000000",
        479 => "00000000",
        480 => "00000000",
        481 => "00000000",
        482 => "01001000",
        483 => "11011011",
        484 => "01001000",
        485 => "00000000",
        486 => "00000000",
        487 => "01001000",
        488 => "11011011",
        489 => "01001000",
        490 => "00000000",
        491 => "00000000",
        492 => "00000000",
        493 => "00000000",
        494 => "00000000",
        495 => "11011010",
        496 => "11011010",
        497 => "00000000",
        498 => "00000000",
        499 => "10110110",
        500 => "11011010",
        501 => "00000000",
        502 => "00000000",
        503 => "00000000",
        504 => "00000000",
        505 => "00000000",
        506 => "00000000",
        507 => "00000000",
        508 => "11011010",
        509 => "11111111",
        510 => "11111111",
        511 => "11011011",
        512 => "00100100",
        513 => "00000000",
        514 => "00000000",
        515 => "00000000",
        516 => "00000000",
        517 => "00000000",
        518 => "00000000",
        519 => "00000000",
        520 => "00000000",
        521 => "00000000",
        522 => "00000000",
        523 => "00000000",
        524 => "00000000",
        525 => "00000000",
        526 => "00000000",
        527 => "00000000",
        528 => "00000000",
        529 => "00000000",
        530 => "00000000",
        531 => "00000000",
        532 => "00000000",
        533 => "00000000",
        534 => "00000000",
        535 => "00000000",
        536 => "00000000",
        537 => "00000000",
        538 => "00000000",
        539 => "00000000",
        540 => "00000000",
        541 => "00000000",
        542 => "00000000",
        543 => "10110110",
        544 => "11111111",
        545 => "11111111",
        546 => "11111111",
        547 => "11111111",
        548 => "11111111",
        549 => "01001000",
        550 => "00000000",
        551 => "00000000",
        552 => "00000000",
        553 => "00000000",
        554 => "01001000",
        555 => "11011011",
        556 => "01001000",
        557 => "00000000",
        558 => "00000000",
        559 => "00000000",
        560 => "00000000",
        561 => "00000000",
        562 => "00000000",
        563 => "00000000",
        564 => "00000000",
        565 => "00000000",
        566 => "01001000",
        567 => "11011011",
        568 => "01001000",
        569 => "00000000",
        570 => "00000000",
        571 => "00000000",
        572 => "00000000",
        573 => "00000000",
        574 => "00000000",
        575 => "00000000",
        576 => "00000000",
        577 => "00000000",
        578 => "00000000",
        579 => "10110110",
        580 => "10110110",
        581 => "00000000",
        582 => "00000000",
        583 => "00000000",
        584 => "00000000",
        585 => "00000000",
        586 => "00000000",
        587 => "00000000",
        588 => "00000000",
        589 => "00000000",
        590 => "00100100",
        591 => "11011011",
        592 => "11111111",
        593 => "11111111",
        594 => "11111111",
        595 => "11111111",
        596 => "11111111",
        597 => "01001000",
        598 => "00000000",
        599 => "00000000",
        600 => "00000000",
        601 => "00000000",
        602 => "00000000",
        603 => "00000000",
        604 => "00000000",
        605 => "00000000",
        606 => "00000000",
        607 => "00000000",
        608 => "00000000",
        609 => "00000000",
        610 => "00000000",
        611 => "00000000",
        612 => "00000000",
        613 => "00000000",
        614 => "00000000",
        615 => "01101101",
        616 => "11111111",
        617 => "11111111",
        618 => "10010001",
        619 => "01001000",
        620 => "11011010",
        621 => "00100100",
        622 => "00000000",
        623 => "00000000",
        624 => "00000000",
        625 => "00000000",
        626 => "00100100",
        627 => "11011010",
        628 => "01101101",
        629 => "10110110",
        630 => "10010001",
        631 => "00100100",
        632 => "11011010",
        633 => "01001000",
        634 => "00000000",
        635 => "00000000",
        636 => "00000000",
        637 => "00000000",
        638 => "01001000",
        639 => "11011010",
        640 => "00100100",
        641 => "10110110",
        642 => "10010001",
        643 => "00100100",
        644 => "11011010",
        645 => "01001000",
        646 => "00000000",
        647 => "00000000",
        648 => "00000000",
        649 => "00000000",
        650 => "00100100",
        651 => "11011011",
        652 => "10010001",
        653 => "10110110",
        654 => "10010001",
        655 => "10010001",
        656 => "11011011",
        657 => "00100100",
        658 => "00000000",
        659 => "00000000",
        660 => "00000000",
        661 => "00000000",
        662 => "00000000",
        663 => "00100100",
        664 => "11011011",
        665 => "11111111",
        666 => "11111111",
        667 => "11111111",
        668 => "01001000",
        669 => "00000000",
        670 => "00000000",
        671 => "00000000",
        672 => "00000000",
        673 => "00000000",
        674 => "00000000",
        675 => "00000000",
        676 => "00000000",
        677 => "00000000",
        678 => "00000000",
        679 => "00000000",
        680 => "00000000",
        681 => "00000000",
        682 => "00000000",
        683 => "00000000",
        684 => "00000000",
        685 => "00000000",
        686 => "00000000",
        687 => "00000000",
        688 => "00000000",
        689 => "00000000",
        690 => "00000000",
        691 => "00000000",
        692 => "00000000",
        693 => "00000000",
        694 => "00000000",
        695 => "00000000",
        696 => "00000000",
        697 => "00000000",
        698 => "00100100",
        699 => "11011011",
        700 => "11111111",
        701 => "11111111",
        702 => "11111111",
        703 => "11111111",
        704 => "11111111",
        705 => "01001000",
        706 => "00000000",
        707 => "00000000",
        708 => "00000000",
        709 => "00000000",
        710 => "00000000",
        711 => "00000000",
        712 => "00000000",
        713 => "00000000",
        714 => "00000000",
        715 => "10110110",
        716 => "10110110",
        717 => "00000000",
        718 => "00000000",
        719 => "00000000",
        720 => "00000000",
        721 => "00000000",
        722 => "00000000",
        723 => "00000000",
        724 => "00000000",
        725 => "00000000",
        726 => "00000000",
        727 => "00100100",
        728 => "11011010",
        729 => "01001000",
        730 => "00000000",
        731 => "00000000",
        732 => "00000000",
        733 => "00000000",
        734 => "00000000",
        735 => "00000000",
        736 => "00000000",
        737 => "00000000",
        738 => "00000000",
        739 => "01001000",
        740 => "11011011",
        741 => "01001000",
        742 => "00000000",
        743 => "00000000",
        744 => "00000000",
        745 => "00000000",
        746 => "00100100",
        747 => "11011011",
        748 => "11111111",
        749 => "11111111",
        750 => "11111111",
        751 => "11111111",
        752 => "10110110",
        753 => "00000000",
        754 => "00000000",
        755 => "00000000",
        756 => "00000000",
        757 => "00000000",
        758 => "00000000",
        759 => "00000000",
        760 => "00000000",
        761 => "00000000",
        762 => "00000000",
        763 => "00000000",
        764 => "00000000",
        765 => "00000000",
        766 => "00000000",
        767 => "00000000",
        768 => "00000000",
        769 => "00000000",
        770 => "00000000",
        771 => "00000000",
        772 => "00000000",
        773 => "00000000",
        774 => "00000000",
        775 => "00000000",
        776 => "00000000",
        777 => "00000000",
        778 => "00000000",
        779 => "00000000",
        780 => "00000000",
        781 => "00000000",
        782 => "00100100",
        783 => "11011011",
        784 => "11111111",
        785 => "11111111",
        786 => "11111111",
        787 => "11111111",
        788 => "11111111",
        789 => "11111111",
        790 => "11111111",
        791 => "10110110",
        792 => "00000000",
        793 => "00000000",
        794 => "01001000",
        795 => "11011010",
        796 => "00100100",
        797 => "00000000",
        798 => "00000000",
        799 => "11011010",
        800 => "10110110",
        801 => "00000000",
        802 => "00000000",
        803 => "00000000",
        804 => "00000000",
        805 => "00000000",
        806 => "01001000",
        807 => "11011010",
        808 => "00100100",
        809 => "00000000",
        810 => "00000000",
        811 => "00100100",
        812 => "11011010",
        813 => "01001000",
        814 => "00000000",
        815 => "00000000",
        816 => "00000000",
        817 => "00000000",
        818 => "00000000",
        819 => "11011010",
        820 => "10010001",
        821 => "00000000",
        822 => "00000000",
        823 => "01101101",
        824 => "11011011",
        825 => "01001000",
        826 => "00000000",
        827 => "00000000",
        828 => "00000000",
        829 => "00000000",
        830 => "00000000",
        831 => "00100100",
        832 => "11011011",
        833 => "11111111",
        834 => "11111111",
        835 => "11111111",
        836 => "01101101",
        837 => "00000000",
        838 => "00000000",
        839 => "00000000",
        840 => "00000000",
        841 => "00000000",
        842 => "00000000",
        843 => "00000000",
        844 => "00000000",
        845 => "00000000",
        846 => "00000000",
        847 => "00000000",
        848 => "00000000",
        849 => "00000000",
        850 => "00000000",
        851 => "00000000",
        852 => "00000000",
        853 => "00000000",
        854 => "00000000",
        855 => "01101101",
        856 => "11111111",
        857 => "11111111",
        858 => "10010001",
        859 => "01001000",
        860 => "11011010",
        861 => "00100100",
        862 => "00000000",
        863 => "00000000",
        864 => "00000000",
        865 => "00000000",
        866 => "00100100",
        867 => "11011010",
        868 => "01101101",
        869 => "10110110",
        870 => "10010001",
        871 => "00100100",
        872 => "11011010",
        873 => "01001000",
        874 => "00000000",
        875 => "00000000",
        876 => "00000000",
        877 => "00000000",
        878 => "01001000",
        879 => "11011010",
        880 => "00100100",
        881 => "10110110",
        882 => "10010001",
        883 => "00100100",
        884 => "11011010",
        885 => "01001000",
        886 => "00000000",
        887 => "00000000",
        888 => "00000000",
        889 => "00000000",
        890 => "00100100",
        891 => "11011011",
        892 => "10010001",
        893 => "10110110",
        894 => "10010001",
        895 => "10010001",
        896 => "11011011",
        897 => "00100100",
        898 => "00000000",
        899 => "00000000",
        900 => "00000000",
        901 => "00000000",
        902 => "00000000",
        903 => "00100100",
        904 => "11011011",
        905 => "11111111",
        906 => "11111111",
        907 => "11111111",
        908 => "01001000",
        909 => "00000000",
        910 => "00000000",
        911 => "00000000",
        912 => "00000000",
        913 => "00000000",
        914 => "00000000",
        915 => "00000000",
        916 => "00000000",
        917 => "00000000",
        918 => "00000000",
        919 => "00000000",
        920 => "00000000",
        921 => "00000000",
        922 => "00000000",
        923 => "00000000",
        924 => "00000000",
        925 => "00000000",
        926 => "00000000",
        927 => "00000000",
        928 => "00000000",
        929 => "00000000",
        930 => "00000000",
        931 => "00000000",
        932 => "00000000",
        933 => "00000000",
        934 => "00000000",
        935 => "00000000",
        936 => "00000000",
        937 => "00000000",
        938 => "00000000",
        939 => "10110110",
        940 => "11111111",
        941 => "10010001",
        942 => "00000000",
        943 => "00000000",
        944 => "00000000",
        945 => "00000000",
        946 => "00000000",
        947 => "00000000",
        948 => "00000000",
        949 => "00000000",
        950 => "01001000",
        951 => "11011011",
        952 => "01001000",
        953 => "00000000",
        954 => "00000000",
        955 => "00000000",
        956 => "00000000",
        957 => "00000000",
        958 => "00000000",
        959 => "00000000",
        960 => "00000000",
        961 => "00000000",
        962 => "00100100",
        963 => "11011010",
        964 => "01001000",
        965 => "00000000",
        966 => "00000000",
        967 => "00000000",
        968 => "00000000",
        969 => "00000000",
        970 => "00000000",
        971 => "00000000",
        972 => "00000000",
        973 => "00000000",
        974 => "00000000",
        975 => "10010001",
        976 => "11011010",
        977 => "00000000",
        978 => "00000000",
        979 => "00000000",
        980 => "00000000",
        981 => "00000000",
        982 => "00000000",
        983 => "00000000",
        984 => "00000000",
        985 => "00000000",
        986 => "00100100",
        987 => "11011011",
        988 => "11111111",
        989 => "11111111",
        990 => "11111111",
        991 => "11111111",
        992 => "11111111",
        993 => "01001000",
        994 => "00000000",
        995 => "00000000",
        996 => "00000000",
        997 => "00000000",
        998 => "00000000",
        999 => "00000000",
        1000 => "00000000",
        1001 => "00000000",
        1002 => "00000000",
        1003 => "00000000",
        1004 => "00000000",
        1005 => "00000000",
        1006 => "00000000",
        1007 => "00000000",
        1008 => "00000000",
        1009 => "00000000",
        1010 => "00000000",
        1011 => "00000000",
        1012 => "00000000",
        1013 => "00000000",
        1014 => "00000000",
        1015 => "00000000",
        1016 => "00000000",
        1017 => "00000000",
        1018 => "00000000",
        1019 => "00000000",
        1020 => "00000000",
        1021 => "10110110",
        1022 => "01101101",
        1023 => "00000000",
        1024 => "10010001",
        1025 => "10110110",
        1026 => "00000000",
        1027 => "00000000",
        1028 => "00000000",
        1029 => "00000000",
        1030 => "00000000",
        1031 => "00000000",
        1032 => "00000000",
        1033 => "10110110",
        1034 => "01101101",
        1035 => "00000000",
        1036 => "10010001",
        1037 => "10110110",
        1038 => "00000000",
        1039 => "00000000",
        1040 => "00000000",
        1041 => "00000000",
        1042 => "00000000",
        1043 => "00000000",
        1044 => "00000000",
        1045 => "10110110",
        1046 => "01101101",
        1047 => "00000000",
        1048 => "10010001",
        1049 => "10110110",
        1050 => "00000000",
        1051 => "00000000",
        1052 => "00000000",
        1053 => "00000000",
        1054 => "00000000",
        1055 => "00000000",
        1056 => "00000000",
        1057 => "11011010",
        1058 => "11111111",
        1059 => "11111111",
        1060 => "11111111",
        1061 => "11111111",
        1062 => "11111111",
        1063 => "11111111",
        1064 => "11111111",
        1065 => "01001000",
        1066 => "00000000",
        1067 => "00000000");

begin

    process(clk)
    begin
    
        if rising_edge(clk) then
            if rst = '1' then
                Freq <= (others => (others => '0'));
            else
                dout <= Freq(to_integer(unsigned(addr)));
            end if;
        end if;
    end process;


end Behavioral;

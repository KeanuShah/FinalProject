

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity RedClass is
    port(clk: in std_logic;
         addr: in std_logic_vector(11 downto 0);
         dout: out std_logic_vector(7 downto 0));
end RedClass;

architecture Behavioral of RedClass is

    type mem is array (0 to 2623) of std_logic_vector(7 downto 0);
    signal Red: mem := (
        0 => "00000001",
1 => "00000001",
2 => "00000001",
3 => "00000001",
4 => "00000001",
5 => "00000001",
6 => "00000001",
7 => "00000001",
8 => "00000001",
9 => "00000001",
10 => "00000001",
11 => "00000001",
12 => "00000001",
13 => "00000001",
14 => "00000001",
15 => "00000001",
16 => "00000001",
17 => "00000001",
18 => "00000001",
19 => "00000001",
20 => "00000001",
21 => "00000001",
22 => "00000001",
23 => "00000001",
24 => "00000001",
25 => "00000001",
26 => "00000001",
27 => "00000001",
28 => "00000001",
29 => "00000001",
30 => "00000001",
31 => "00000001",
32 => "00000001",
33 => "00000001",
34 => "00000001",
35 => "00000001",
36 => "00000001",
37 => "00000001",
38 => "00000001",
39 => "00000001",
40 => "00000001",
41 => "00000001",
42 => "00000001",
43 => "00000001",
44 => "00000001",
45 => "00000001",
46 => "00000001",
47 => "00000001",
48 => "00000001",
49 => "00000001",
50 => "00000001",
51 => "00000001",
52 => "00000001",
53 => "00000001",
54 => "00000001",
55 => "00000001",
56 => "00000001",
57 => "00000001",
58 => "00000001",
59 => "00000001",
60 => "00000001",
61 => "00000001",
62 => "00000001",
63 => "00000001",
64 => "00000001",
65 => "00000001",
66 => "00000001",
67 => "00000001",
68 => "00000001",
69 => "00000001",
70 => "00000001",
71 => "00000001",
72 => "00000001",
73 => "00000001",
74 => "00000001",
75 => "00000001",
76 => "00000001",
77 => "00000001",
78 => "00000001",
79 => "00000001",
80 => "00000001",
81 => "00000001",
82 => "00000001",
83 => "00000001",
84 => "00100101",
85 => "10110110",
86 => "11111111",
87 => "11111111",
88 => "11111111",
89 => "11111111",
90 => "11111111",
91 => "11111111",
92 => "11111111",
93 => "11111111",
94 => "11111111",
95 => "11111111",
96 => "11111111",
97 => "11111111",
98 => "11111111",
99 => "11111111",
100 => "11111111",
101 => "11111111",
102 => "11111111",
103 => "11111111",
104 => "11111111",
105 => "11111111",
106 => "11111111",
107 => "11111111",
108 => "11111111",
109 => "11111111",
110 => "11111111",
111 => "11111111",
112 => "11111111",
113 => "11111111",
114 => "11111111",
115 => "11111111",
116 => "11111111",
117 => "11111111",
118 => "11111111",
119 => "11111111",
120 => "11111111",
121 => "11111111",
122 => "11111111",
123 => "11111111",
124 => "11111111",
125 => "11111111",
126 => "11111111",
127 => "11111111",
128 => "11111111",
129 => "11111111",
130 => "11111111",
131 => "11111111",
132 => "11111111",
133 => "11111111",
134 => "11111111",
135 => "11111111",
136 => "11111111",
137 => "11111111",
138 => "11111111",
139 => "11111111",
140 => "11111111",
141 => "11111111",
142 => "11111111",
143 => "11111111",
144 => "11111111",
145 => "11111111",
146 => "11111111",
147 => "11111111",
148 => "11111111",
149 => "11111111",
150 => "11111111",
151 => "11111111",
152 => "11111111",
153 => "11111111",
154 => "11111111",
155 => "11111111",
156 => "11111111",
157 => "11111111",
158 => "11111111",
159 => "11111111",
160 => "10110110",
161 => "00100101",
162 => "00000001",
163 => "00000001",
164 => "00000001",
165 => "00100101",
166 => "11111111",
167 => "10101001",
168 => "10000000",
169 => "10000000",
170 => "10000000",
171 => "10000000",
172 => "10000000",
173 => "10000000",
174 => "10000000",
175 => "10000000",
176 => "10000000",
177 => "10000000",
178 => "10000000",
179 => "10000000",
180 => "10000000",
181 => "10000000",
182 => "10000000",
183 => "10000000",
184 => "10000000",
185 => "10000000",
186 => "10000000",
187 => "10000000",
188 => "10000000",
189 => "10000000",
190 => "10000000",
191 => "10000000",
192 => "10000000",
193 => "10000000",
194 => "10000000",
195 => "10000000",
196 => "10000000",
197 => "10000000",
198 => "10000000",
199 => "10000000",
200 => "10000000",
201 => "10000000",
202 => "10000000",
203 => "10000000",
204 => "10000000",
205 => "10000000",
206 => "10000000",
207 => "10000000",
208 => "10000000",
209 => "10000000",
210 => "10000000",
211 => "10000000",
212 => "10000000",
213 => "10000000",
214 => "10000000",
215 => "10000000",
216 => "10000000",
217 => "10000000",
218 => "10000000",
219 => "10000000",
220 => "10000000",
221 => "10000000",
222 => "10000000",
223 => "10000000",
224 => "10000000",
225 => "10000000",
226 => "10000000",
227 => "10000000",
228 => "10000000",
229 => "10000000",
230 => "10000000",
231 => "10000000",
232 => "10000000",
233 => "10000000",
234 => "10000000",
235 => "10000000",
236 => "10000000",
237 => "10000000",
238 => "10000000",
239 => "10000000",
240 => "10000000",
241 => "10000000",
242 => "10101001",
243 => "11111111",
244 => "00100101",
245 => "00000001",
246 => "00000001",
247 => "10110110",
248 => "10101001",
249 => "10000000",
250 => "10000000",
251 => "10000000",
252 => "10000000",
253 => "10000000",
254 => "10000000",
255 => "10000000",
256 => "10000000",
257 => "10000000",
258 => "10000000",
259 => "10000000",
260 => "10000000",
261 => "10000000",
262 => "10000000",
263 => "10000000",
264 => "10000000",
265 => "10000000",
266 => "10000000",
267 => "10000000",
268 => "10000000",
269 => "10000000",
270 => "10000000",
271 => "10000000",
272 => "10000000",
273 => "10000000",
274 => "10000000",
275 => "10000000",
276 => "10000000",
277 => "10000000",
278 => "10000000",
279 => "10000000",
280 => "10000000",
281 => "10000000",
282 => "10000000",
283 => "10000000",
284 => "10000000",
285 => "10000000",
286 => "10000000",
287 => "10000000",
288 => "10000000",
289 => "10000000",
290 => "10000000",
291 => "10000000",
292 => "10000000",
293 => "10000000",
294 => "10000000",
295 => "10000000",
296 => "10000000",
297 => "10000000",
298 => "10000000",
299 => "10000000",
300 => "10000000",
301 => "10000000",
302 => "10000000",
303 => "10000000",
304 => "10000000",
305 => "10000000",
306 => "10000000",
307 => "10000000",
308 => "10000000",
309 => "10000000",
310 => "10000000",
311 => "10000000",
312 => "10000000",
313 => "10000000",
314 => "10000000",
315 => "10000000",
316 => "10000000",
317 => "10000000",
318 => "10000000",
319 => "10000000",
320 => "10000000",
321 => "10000000",
322 => "10000000",
323 => "10000000",
324 => "10000000",
325 => "10101001",
326 => "10110110",
327 => "00000001",
328 => "00000001",
329 => "11111111",
330 => "10000000",
331 => "10000000",
332 => "10000000",
333 => "10000000",
334 => "10000000",
335 => "10000000",
336 => "10000000",
337 => "10000000",
338 => "10000000",
339 => "10000000",
340 => "10000000",
341 => "10000000",
342 => "10000000",
343 => "10000000",
344 => "10000000",
345 => "10000000",
346 => "10000000",
347 => "10000000",
348 => "10000000",
349 => "10000000",
350 => "10000000",
351 => "10000000",
352 => "10000000",
353 => "10000000",
354 => "10000000",
355 => "10000000",
356 => "10000000",
357 => "10000000",
358 => "10000000",
359 => "10000000",
360 => "10000000",
361 => "10000000",
362 => "10000000",
363 => "10000000",
364 => "10000000",
365 => "10000000",
366 => "10000000",
367 => "10000000",
368 => "10000000",
369 => "10000000",
370 => "10000000",
371 => "10000000",
372 => "10000000",
373 => "10000000",
374 => "10000000",
375 => "10000000",
376 => "10000000",
377 => "10000000",
378 => "10000000",
379 => "10000000",
380 => "10000000",
381 => "10000000",
382 => "10000000",
383 => "10000000",
384 => "10000000",
385 => "10000000",
386 => "10000000",
387 => "10000000",
388 => "10000000",
389 => "10000000",
390 => "10000000",
391 => "10000000",
392 => "10000000",
393 => "10000000",
394 => "10000000",
395 => "10000000",
396 => "10000000",
397 => "10000000",
398 => "10000000",
399 => "10000000",
400 => "10000000",
401 => "10000000",
402 => "10000000",
403 => "10000000",
404 => "10000000",
405 => "10000000",
406 => "10000000",
407 => "10000000",
408 => "11111111",
409 => "00000001",
410 => "00000001",
411 => "11111111",
412 => "10000000",
413 => "10000000",
414 => "10000000",
415 => "10000000",
416 => "10000000",
417 => "10000000",
418 => "10000000",
419 => "10000000",
420 => "10000000",
421 => "10000000",
422 => "10000000",
423 => "10000000",
424 => "10000000",
425 => "10000000",
426 => "10000000",
427 => "10000000",
428 => "10000000",
429 => "10000000",
430 => "10000000",
431 => "10000000",
432 => "10000000",
433 => "10000000",
434 => "10000000",
435 => "10000000",
436 => "10000000",
437 => "10000000",
438 => "10000000",
439 => "10000000",
440 => "10000000",
441 => "10000000",
442 => "10000000",
443 => "10000000",
444 => "10000000",
445 => "10000000",
446 => "10000000",
447 => "10000000",
448 => "10000000",
449 => "10000000",
450 => "10000000",
451 => "10000000",
452 => "10000000",
453 => "10000000",
454 => "10000000",
455 => "10000000",
456 => "10000000",
457 => "10000000",
458 => "10000000",
459 => "10000000",
460 => "10000000",
461 => "10000000",
462 => "10000000",
463 => "10000000",
464 => "10000000",
465 => "10000000",
466 => "10000000",
467 => "10000000",
468 => "10000000",
469 => "10000000",
470 => "10000000",
471 => "10000000",
472 => "10000000",
473 => "10000000",
474 => "10000000",
475 => "10000000",
476 => "10000000",
477 => "10000000",
478 => "10000000",
479 => "10000000",
480 => "10000000",
481 => "10000000",
482 => "10000000",
483 => "10000000",
484 => "10000000",
485 => "10000000",
486 => "10000000",
487 => "10000000",
488 => "10000000",
489 => "10000000",
490 => "11111111",
491 => "00000001",
492 => "00000001",
493 => "11111111",
494 => "10000000",
495 => "10000000",
496 => "10000000",
497 => "10000000",
498 => "10000000",
499 => "10000000",
500 => "10000000",
501 => "10000000",
502 => "10000000",
503 => "10000000",
504 => "10000000",
505 => "10000000",
506 => "10000000",
507 => "10000000",
508 => "10000000",
509 => "10000000",
510 => "10000000",
511 => "10000000",
512 => "10000000",
513 => "10000000",
514 => "10000000",
515 => "10000000",
516 => "10000000",
517 => "10000000",
518 => "10000000",
519 => "10000000",
520 => "10000000",
521 => "10000000",
522 => "10000000",
523 => "10000000",
524 => "10000000",
525 => "10000000",
526 => "10000000",
527 => "10000000",
528 => "10000000",
529 => "10000000",
530 => "10000000",
531 => "10000000",
532 => "10000000",
533 => "10000000",
534 => "10000000",
535 => "10000000",
536 => "10000000",
537 => "10000000",
538 => "10000000",
539 => "10000000",
540 => "10000000",
541 => "10000000",
542 => "10000000",
543 => "10000000",
544 => "10000000",
545 => "10000000",
546 => "10000000",
547 => "10000000",
548 => "10000000",
549 => "10000000",
550 => "10000000",
551 => "10000000",
552 => "10000000",
553 => "10000000",
554 => "10000000",
555 => "10000000",
556 => "10000000",
557 => "10000000",
558 => "10000000",
559 => "10000000",
560 => "10000000",
561 => "10000000",
562 => "10000000",
563 => "10000000",
564 => "10000000",
565 => "10000000",
566 => "10000000",
567 => "10000000",
568 => "10000000",
569 => "10000000",
570 => "10000000",
571 => "10000000",
572 => "11111111",
573 => "00000001",
574 => "00000001",
575 => "11111111",
576 => "10000000",
577 => "10000000",
578 => "10000000",
579 => "10000000",
580 => "10000000",
581 => "10000000",
582 => "10000000",
583 => "10000000",
584 => "10000000",
585 => "10000000",
586 => "10000000",
587 => "10000000",
588 => "10000000",
589 => "10000000",
590 => "10000000",
591 => "10000000",
592 => "10000000",
593 => "10000000",
594 => "10000000",
595 => "10000000",
596 => "10000000",
597 => "10000000",
598 => "10000000",
599 => "10000000",
600 => "10000000",
601 => "10000000",
602 => "10000000",
603 => "10000000",
604 => "10000000",
605 => "10000000",
606 => "10000000",
607 => "10000000",
608 => "10000000",
609 => "10000000",
610 => "10000000",
611 => "10000000",
612 => "10000000",
613 => "10000000",
614 => "10000000",
615 => "10000000",
616 => "10000000",
617 => "10000000",
618 => "10000000",
619 => "10000000",
620 => "10000000",
621 => "10000000",
622 => "10000000",
623 => "10000000",
624 => "10000000",
625 => "10000000",
626 => "10000000",
627 => "10000000",
628 => "10000000",
629 => "10000000",
630 => "10000000",
631 => "10000000",
632 => "10000000",
633 => "10000000",
634 => "10000000",
635 => "10000000",
636 => "10000000",
637 => "10000000",
638 => "10000000",
639 => "10000000",
640 => "10000000",
641 => "10000000",
642 => "10000000",
643 => "10000000",
644 => "10000000",
645 => "10000000",
646 => "10000000",
647 => "10000000",
648 => "10000000",
649 => "10000000",
650 => "10000000",
651 => "10000000",
652 => "10000000",
653 => "10000000",
654 => "11111111",
655 => "00000001",
656 => "00000001",
657 => "11111111",
658 => "10000000",
659 => "10000000",
660 => "10000000",
661 => "10000000",
662 => "10000000",
663 => "10000000",
664 => "10000000",
665 => "10000000",
666 => "10000000",
667 => "10000000",
668 => "10000000",
669 => "10000000",
670 => "10000000",
671 => "10000000",
672 => "10000000",
673 => "10000000",
674 => "10000000",
675 => "10000000",
676 => "10000000",
677 => "10000000",
678 => "10000000",
679 => "10000000",
680 => "10000000",
681 => "10000000",
682 => "10000000",
683 => "10000000",
684 => "10000000",
685 => "10000000",
686 => "10000000",
687 => "10000000",
688 => "10000000",
689 => "10000000",
690 => "10000000",
691 => "10000000",
692 => "10000000",
693 => "10000000",
694 => "10000000",
695 => "10000000",
696 => "10000000",
697 => "10000000",
698 => "10000000",
699 => "10000000",
700 => "10000000",
701 => "10000000",
702 => "10000000",
703 => "10000000",
704 => "10000000",
705 => "10000000",
706 => "10000000",
707 => "10000000",
708 => "10000000",
709 => "10000000",
710 => "10000000",
711 => "10000000",
712 => "10000000",
713 => "10000000",
714 => "10000000",
715 => "10000000",
716 => "10000000",
717 => "10000000",
718 => "10000000",
719 => "10000000",
720 => "10000000",
721 => "10000000",
722 => "10000000",
723 => "10000000",
724 => "10000000",
725 => "10000000",
726 => "10000000",
727 => "10000000",
728 => "10000000",
729 => "10000000",
730 => "10000000",
731 => "10000000",
732 => "10000000",
733 => "10000000",
734 => "10000000",
735 => "10000000",
736 => "11111111",
737 => "00000001",
738 => "00000001",
739 => "11111111",
740 => "10000000",
741 => "10000000",
742 => "10000000",
743 => "10000000",
744 => "10000000",
745 => "10000000",
746 => "10000000",
747 => "10000000",
748 => "10000000",
749 => "10000000",
750 => "10000000",
751 => "10000000",
752 => "10000000",
753 => "10000000",
754 => "10000000",
755 => "10000000",
756 => "10000000",
757 => "10000000",
758 => "10000000",
759 => "10000000",
760 => "10000000",
761 => "10000000",
762 => "10000000",
763 => "10000000",
764 => "10000000",
765 => "10000000",
766 => "10000000",
767 => "10000000",
768 => "10000000",
769 => "10000000",
770 => "10000000",
771 => "10000000",
772 => "10000000",
773 => "10000000",
774 => "10000000",
775 => "10000000",
776 => "10000000",
777 => "10000000",
778 => "10000000",
779 => "10000000",
780 => "10000000",
781 => "10000000",
782 => "10000000",
783 => "10000000",
784 => "10000000",
785 => "10000000",
786 => "10000000",
787 => "10000000",
788 => "10000000",
789 => "10000000",
790 => "10000000",
791 => "10000000",
792 => "10000000",
793 => "10000000",
794 => "10000000",
795 => "10000000",
796 => "10000000",
797 => "10000000",
798 => "10000000",
799 => "10000000",
800 => "10000000",
801 => "10000000",
802 => "10000000",
803 => "10000000",
804 => "10000000",
805 => "10000000",
806 => "10000000",
807 => "10000000",
808 => "10000000",
809 => "10000000",
810 => "10000000",
811 => "10000000",
812 => "10000000",
813 => "10000000",
814 => "10000000",
815 => "10000000",
816 => "10000000",
817 => "10000000",
818 => "11111111",
819 => "00000001",
820 => "00000001",
821 => "11111111",
822 => "10000000",
823 => "10000000",
824 => "10000000",
825 => "10000000",
826 => "10000000",
827 => "10000000",
828 => "10000000",
829 => "10000000",
830 => "10000000",
831 => "10000000",
832 => "10000000",
833 => "10000000",
834 => "10000000",
835 => "10000000",
836 => "10000000",
837 => "10000000",
838 => "10000000",
839 => "10000000",
840 => "10000000",
841 => "10000000",
842 => "10000000",
843 => "10000000",
844 => "10000000",
845 => "10000000",
846 => "10000000",
847 => "10000000",
848 => "10000000",
849 => "10000000",
850 => "10000000",
851 => "10000000",
852 => "10000000",
853 => "10000000",
854 => "10000000",
855 => "10000000",
856 => "10000000",
857 => "10000000",
858 => "10000000",
859 => "10000000",
860 => "10000000",
861 => "10000000",
862 => "10000000",
863 => "10000000",
864 => "10000000",
865 => "10000000",
866 => "10000000",
867 => "10000000",
868 => "10000000",
869 => "10000000",
870 => "10000000",
871 => "10000000",
872 => "10000000",
873 => "10000000",
874 => "10000000",
875 => "10000000",
876 => "10000000",
877 => "10000000",
878 => "10000000",
879 => "10000000",
880 => "10000000",
881 => "10000000",
882 => "10000000",
883 => "10000000",
884 => "10000000",
885 => "10000000",
886 => "10000000",
887 => "10000000",
888 => "10000000",
889 => "10000000",
890 => "10000000",
891 => "10000000",
892 => "10000000",
893 => "10000000",
894 => "10000000",
895 => "10000000",
896 => "10000000",
897 => "10000000",
898 => "10000000",
899 => "10000000",
900 => "11111111",
901 => "00000001",
902 => "00000001",
903 => "11111111",
904 => "10000000",
905 => "10000000",
906 => "10000000",
907 => "10000000",
908 => "10000000",
909 => "10000000",
910 => "10000000",
911 => "10000000",
912 => "10000000",
913 => "10000000",
914 => "10000000",
915 => "10000000",
916 => "10000000",
917 => "10000000",
918 => "10000000",
919 => "10000000",
920 => "10000000",
921 => "10000000",
922 => "10000000",
923 => "10000000",
924 => "10000000",
925 => "10000000",
926 => "10000000",
927 => "10000000",
928 => "10000000",
929 => "10000000",
930 => "10000000",
931 => "10000000",
932 => "10000000",
933 => "10000000",
934 => "10000000",
935 => "10000000",
936 => "10000000",
937 => "10000000",
938 => "10000000",
939 => "10000000",
940 => "10000000",
941 => "10000000",
942 => "10000000",
943 => "10000000",
944 => "10000000",
945 => "10000000",
946 => "10000000",
947 => "10000000",
948 => "10000000",
949 => "10000000",
950 => "10000000",
951 => "10000000",
952 => "10000000",
953 => "10000000",
954 => "10000000",
955 => "10000000",
956 => "10000000",
957 => "10000000",
958 => "10000000",
959 => "10000000",
960 => "10000000",
961 => "10000000",
962 => "10000000",
963 => "10000000",
964 => "10000000",
965 => "10000000",
966 => "10000000",
967 => "10000000",
968 => "10000000",
969 => "10000000",
970 => "10000000",
971 => "10000000",
972 => "10000000",
973 => "10000000",
974 => "10000000",
975 => "10000000",
976 => "10000000",
977 => "10000000",
978 => "10000000",
979 => "10000000",
980 => "10000000",
981 => "10000000",
982 => "11111111",
983 => "00000001",
984 => "00000001",
985 => "11111111",
986 => "10000000",
987 => "10000000",
988 => "10000000",
989 => "10000000",
990 => "10000000",
991 => "10000000",
992 => "10000000",
993 => "10000000",
994 => "10000000",
995 => "10000000",
996 => "10000000",
997 => "10000000",
998 => "10000000",
999 => "10000000",
1000 => "10000000",
1001 => "10000000",
1002 => "10000000",
1003 => "10000000",
1004 => "10000000",
1005 => "10000000",
1006 => "10000001",
1007 => "11011011",
1008 => "11111111",
1009 => "11111111",
1010 => "11111110",
1011 => "11000000",
1012 => "10000000",
1013 => "10000000",
1014 => "10000000",
1015 => "10000000",
1016 => "10000000",
1017 => "10000000",
1018 => "10000000",
1019 => "10000000",
1020 => "10000000",
1021 => "10000000",
1022 => "10000000",
1023 => "10000000",
1024 => "10000000",
1025 => "10000000",
1026 => "10000000",
1027 => "10000000",
1028 => "10000000",
1029 => "10000000",
1030 => "10000000",
1031 => "10000000",
1032 => "10000000",
1033 => "10000000",
1034 => "10000000",
1035 => "10000000",
1036 => "10000000",
1037 => "10000000",
1038 => "10000000",
1039 => "10000000",
1040 => "10000000",
1041 => "10000000",
1042 => "10000000",
1043 => "10000000",
1044 => "10000000",
1045 => "10000000",
1046 => "10000000",
1047 => "10000000",
1048 => "10000000",
1049 => "10000000",
1050 => "10000000",
1051 => "10000000",
1052 => "10000000",
1053 => "10000000",
1054 => "10000000",
1055 => "10000000",
1056 => "10000000",
1057 => "10000000",
1058 => "10000000",
1059 => "10000000",
1060 => "10000000",
1061 => "10000000",
1062 => "10000000",
1063 => "10000000",
1064 => "11111111",
1065 => "00000001",
1066 => "00000001",
1067 => "11111111",
1068 => "10000000",
1069 => "10000000",
1070 => "10000000",
1071 => "10000000",
1072 => "10000000",
1073 => "10000000",
1074 => "10000000",
1075 => "10000000",
1076 => "10000000",
1077 => "10000000",
1078 => "10000000",
1079 => "10000000",
1080 => "10000000",
1081 => "10000000",
1082 => "10000000",
1083 => "10000000",
1084 => "10000000",
1085 => "10000000",
1086 => "10000000",
1087 => "10000000",
1088 => "11011011",
1089 => "11111010",
1090 => "11000000",
1091 => "10000000",
1092 => "10000000",
1093 => "10000000",
1094 => "10000000",
1095 => "10000000",
1096 => "10000000",
1097 => "10000000",
1098 => "10000000",
1099 => "10000000",
1100 => "10000000",
1101 => "10000000",
1102 => "10000000",
1103 => "10000000",
1104 => "10000000",
1105 => "10000000",
1106 => "10000000",
1107 => "10000000",
1108 => "10000000",
1109 => "10000000",
1110 => "10000000",
1111 => "10000000",
1112 => "10000000",
1113 => "10000000",
1114 => "10000000",
1115 => "10000000",
1116 => "10000000",
1117 => "10000000",
1118 => "10000000",
1119 => "10000000",
1120 => "10000000",
1121 => "10000000",
1122 => "10000000",
1123 => "10000000",
1124 => "10000000",
1125 => "10000000",
1126 => "10000000",
1127 => "10000000",
1128 => "10000000",
1129 => "10000000",
1130 => "10000000",
1131 => "10000000",
1132 => "10000000",
1133 => "10000000",
1134 => "10000000",
1135 => "10000000",
1136 => "10000000",
1137 => "10000000",
1138 => "10000000",
1139 => "10000000",
1140 => "10000000",
1141 => "10000000",
1142 => "10000000",
1143 => "10000000",
1144 => "10000000",
1145 => "10000000",
1146 => "11111111",
1147 => "00000001",
1148 => "00000001",
1149 => "11111111",
1150 => "10000000",
1151 => "10000000",
1152 => "10000000",
1153 => "10000000",
1154 => "10000000",
1155 => "10000000",
1156 => "10000000",
1157 => "10000000",
1158 => "10000000",
1159 => "10000000",
1160 => "10000000",
1161 => "10000000",
1162 => "10000000",
1163 => "10000000",
1164 => "10000000",
1165 => "10000000",
1166 => "10000000",
1167 => "10000000",
1168 => "10000000",
1169 => "10000001",
1170 => "11011011",
1171 => "11111010",
1172 => "11000000",
1173 => "10000000",
1174 => "10000000",
1175 => "10000000",
1176 => "10000000",
1177 => "10000001",
1178 => "11011011",
1179 => "11111111",
1180 => "11111111",
1181 => "11110101",
1182 => "10000001",
1183 => "11011011",
1184 => "11111001",
1185 => "10000000",
1186 => "10000000",
1187 => "10010010",
1188 => "11111111",
1189 => "11001100",
1190 => "10000000",
1191 => "11011011",
1192 => "11111111",
1193 => "11111111",
1194 => "11111001",
1195 => "10000000",
1196 => "10000001",
1197 => "11111111",
1198 => "11111010",
1199 => "11111111",
1200 => "11111111",
1201 => "11111001",
1202 => "10000000",
1203 => "10000000",
1204 => "11011011",
1205 => "11111111",
1206 => "11111111",
1207 => "11111001",
1208 => "10000000",
1209 => "10000000",
1210 => "10000000",
1211 => "10000000",
1212 => "10000000",
1213 => "10000000",
1214 => "10000000",
1215 => "10000000",
1216 => "10000000",
1217 => "10000000",
1218 => "10000000",
1219 => "10000000",
1220 => "10000000",
1221 => "10000000",
1222 => "10000000",
1223 => "10000000",
1224 => "10000000",
1225 => "10000000",
1226 => "10000000",
1227 => "10000000",
1228 => "11111111",
1229 => "00000001",
1230 => "00000001",
1231 => "11111111",
1232 => "10000000",
1233 => "10000000",
1234 => "10000000",
1235 => "10000000",
1236 => "10000000",
1237 => "10000000",
1238 => "10000000",
1239 => "10000000",
1240 => "10000000",
1241 => "10000000",
1242 => "10000000",
1243 => "10000000",
1244 => "10000000",
1245 => "10000000",
1246 => "10000000",
1247 => "10000000",
1248 => "10000000",
1249 => "10000000",
1250 => "10000000",
1251 => "10000000",
1252 => "10010010",
1253 => "11111111",
1254 => "11111111",
1255 => "11111110",
1256 => "11000000",
1257 => "10000000",
1258 => "10000000",
1259 => "11011011",
1260 => "11111001",
1261 => "10000000",
1262 => "10001110",
1263 => "11111111",
1264 => "11110000",
1265 => "11010111",
1266 => "11111110",
1267 => "11000000",
1268 => "10000000",
1269 => "11011011",
1270 => "11111001",
1271 => "10000000",
1272 => "11010111",
1273 => "11111010",
1274 => "11000000",
1275 => "10000001",
1276 => "11111111",
1277 => "11110101",
1278 => "10000001",
1279 => "11111111",
1280 => "11111110",
1281 => "11000000",
1282 => "10010010",
1283 => "11111111",
1284 => "11001100",
1285 => "11010111",
1286 => "11111010",
1287 => "11000000",
1288 => "10000001",
1289 => "11111111",
1290 => "11110101",
1291 => "10000000",
1292 => "10000000",
1293 => "10000000",
1294 => "10000000",
1295 => "10000000",
1296 => "10000000",
1297 => "10000000",
1298 => "10000000",
1299 => "10000000",
1300 => "10000000",
1301 => "10000000",
1302 => "10000000",
1303 => "10000000",
1304 => "10000000",
1305 => "10000000",
1306 => "10000000",
1307 => "10000000",
1308 => "10000000",
1309 => "10000000",
1310 => "11111111",
1311 => "00000001",
1312 => "00000001",
1313 => "11111111",
1314 => "10000000",
1315 => "10000000",
1316 => "10000000",
1317 => "10000000",
1318 => "10000000",
1319 => "10000000",
1320 => "10000000",
1321 => "10000000",
1322 => "10000000",
1323 => "10000000",
1324 => "10000000",
1325 => "10000000",
1326 => "10000000",
1327 => "10000000",
1328 => "10000000",
1329 => "10000000",
1330 => "10000000",
1331 => "10000000",
1332 => "10000000",
1333 => "10000000",
1334 => "10000000",
1335 => "10000000",
1336 => "11011011",
1337 => "11111111",
1338 => "11111111",
1339 => "11110000",
1340 => "10000001",
1341 => "11111111",
1342 => "11111111",
1343 => "11111111",
1344 => "11111111",
1345 => "11111111",
1346 => "11110000",
1347 => "10000001",
1348 => "11111111",
1349 => "11110000",
1350 => "10000001",
1351 => "11111111",
1352 => "11110000",
1353 => "10000001",
1354 => "11011011",
1355 => "11111111",
1356 => "11111111",
1357 => "11111111",
1358 => "11111111",
1359 => "11110101",
1360 => "10000001",
1361 => "11111111",
1362 => "11110101",
1363 => "10000000",
1364 => "10000000",
1365 => "10000000",
1366 => "10000001",
1367 => "11011011",
1368 => "11111111",
1369 => "11111111",
1370 => "11111111",
1371 => "11111111",
1372 => "11110101",
1373 => "10000000",
1374 => "10000000",
1375 => "10000000",
1376 => "10000000",
1377 => "10000000",
1378 => "10000000",
1379 => "10000000",
1380 => "10000000",
1381 => "10000000",
1382 => "10000000",
1383 => "10000000",
1384 => "10000000",
1385 => "10000000",
1386 => "10000000",
1387 => "10000000",
1388 => "10000000",
1389 => "10000000",
1390 => "10000000",
1391 => "10000000",
1392 => "11111111",
1393 => "00000001",
1394 => "00000001",
1395 => "11111111",
1396 => "10000000",
1397 => "10000000",
1398 => "10000000",
1399 => "10000000",
1400 => "10000000",
1401 => "10000000",
1402 => "10000000",
1403 => "10000000",
1404 => "10000000",
1405 => "10000000",
1406 => "10000000",
1407 => "10000000",
1408 => "10000000",
1409 => "10000000",
1410 => "10000000",
1411 => "10000000",
1412 => "10000000",
1413 => "10000000",
1414 => "10000000",
1415 => "10000000",
1416 => "10000000",
1417 => "10000000",
1418 => "10000000",
1419 => "10001110",
1420 => "11111111",
1421 => "11110101",
1422 => "10000001",
1423 => "11111111",
1424 => "11110101",
1425 => "10000000",
1426 => "10000000",
1427 => "10000000",
1428 => "10000000",
1429 => "10000000",
1430 => "11011011",
1431 => "11111001",
1432 => "10010010",
1433 => "11111110",
1434 => "11000000",
1435 => "10000001",
1436 => "11011011",
1437 => "11111001",
1438 => "10000000",
1439 => "10000000",
1440 => "10000000",
1441 => "10000000",
1442 => "10000001",
1443 => "11111111",
1444 => "11110101",
1445 => "10000000",
1446 => "10000000",
1447 => "10000000",
1448 => "10000001",
1449 => "11011011",
1450 => "11111001",
1451 => "10000000",
1452 => "10000000",
1453 => "10000000",
1454 => "10000000",
1455 => "10000000",
1456 => "10000000",
1457 => "10000000",
1458 => "10000000",
1459 => "10000000",
1460 => "10000000",
1461 => "10000000",
1462 => "10000000",
1463 => "10000000",
1464 => "10000000",
1465 => "10000000",
1466 => "10000000",
1467 => "10000000",
1468 => "10000000",
1469 => "10000000",
1470 => "10000000",
1471 => "10000000",
1472 => "10000000",
1473 => "10000000",
1474 => "11111111",
1475 => "00000001",
1476 => "00000001",
1477 => "11111111",
1478 => "10000000",
1479 => "10000000",
1480 => "10000000",
1481 => "10000000",
1482 => "10000000",
1483 => "10000000",
1484 => "10000000",
1485 => "10000000",
1486 => "10000000",
1487 => "10000000",
1488 => "10000000",
1489 => "10000000",
1490 => "10000000",
1491 => "10000000",
1492 => "10000000",
1493 => "10000000",
1494 => "10000000",
1495 => "10000000",
1496 => "10000000",
1497 => "10000000",
1498 => "10000000",
1499 => "10000000",
1500 => "10000000",
1501 => "10010010",
1502 => "11111111",
1503 => "11110000",
1504 => "10000001",
1505 => "11011011",
1506 => "11111110",
1507 => "11000000",
1508 => "10000000",
1509 => "10000000",
1510 => "10000000",
1511 => "10000000",
1512 => "10001110",
1513 => "11111110",
1514 => "11111011",
1515 => "11110101",
1516 => "10000000",
1517 => "10000000",
1518 => "11011011",
1519 => "11111111",
1520 => "11001100",
1521 => "10000000",
1522 => "10000000",
1523 => "10000000",
1524 => "10000001",
1525 => "11111111",
1526 => "11110101",
1527 => "10000000",
1528 => "10000000",
1529 => "10000000",
1530 => "10000000",
1531 => "11011011",
1532 => "11111111",
1533 => "11001100",
1534 => "10000000",
1535 => "10000000",
1536 => "10000000",
1537 => "10000000",
1538 => "10000000",
1539 => "10000000",
1540 => "10000000",
1541 => "10000000",
1542 => "10000000",
1543 => "10000000",
1544 => "10000000",
1545 => "10000000",
1546 => "10000000",
1547 => "10000000",
1548 => "10000000",
1549 => "10000000",
1550 => "10000000",
1551 => "10000000",
1552 => "10000000",
1553 => "10000000",
1554 => "10000000",
1555 => "10000000",
1556 => "11111111",
1557 => "00000001",
1558 => "00000001",
1559 => "11111111",
1560 => "10000000",
1561 => "10000000",
1562 => "10000000",
1563 => "10000000",
1564 => "10000000",
1565 => "10000000",
1566 => "10000000",
1567 => "10000000",
1568 => "10000000",
1569 => "10000000",
1570 => "10000000",
1571 => "10000000",
1572 => "10000000",
1573 => "10000000",
1574 => "10000000",
1575 => "10000000",
1576 => "10000000",
1577 => "10000000",
1578 => "10000000",
1579 => "10000001",
1580 => "11011011",
1581 => "11111111",
1582 => "11111111",
1583 => "11111111",
1584 => "11110101",
1585 => "10000000",
1586 => "10000000",
1587 => "10000001",
1588 => "11111111",
1589 => "11111111",
1590 => "11111111",
1591 => "11111111",
1592 => "11001100",
1593 => "10000000",
1594 => "10000001",
1595 => "11011011",
1596 => "11111111",
1597 => "11001100",
1598 => "10000000",
1599 => "10000000",
1600 => "10000001",
1601 => "11011011",
1602 => "11111111",
1603 => "11111111",
1604 => "11111111",
1605 => "11110000",
1606 => "10000001",
1607 => "11111111",
1608 => "11110101",
1609 => "10000000",
1610 => "10000000",
1611 => "10000000",
1612 => "10000000",
1613 => "10000001",
1614 => "11011011",
1615 => "11111111",
1616 => "11111111",
1617 => "11111111",
1618 => "11110000",
1619 => "10000000",
1620 => "10000000",
1621 => "10000000",
1622 => "10000000",
1623 => "10000000",
1624 => "10000000",
1625 => "10000000",
1626 => "10000000",
1627 => "10000000",
1628 => "10000000",
1629 => "10000000",
1630 => "10000000",
1631 => "10000000",
1632 => "10000000",
1633 => "10000000",
1634 => "10000000",
1635 => "10000000",
1636 => "10000000",
1637 => "10000000",
1638 => "11111111",
1639 => "00000001",
1640 => "00000001",
1641 => "11111111",
1642 => "10000000",
1643 => "10000000",
1644 => "10000000",
1645 => "10000000",
1646 => "10000000",
1647 => "10000000",
1648 => "10000000",
1649 => "10000000",
1650 => "10000000",
1651 => "10000000",
1652 => "10000000",
1653 => "10000000",
1654 => "10000000",
1655 => "10000000",
1656 => "10000000",
1657 => "10000000",
1658 => "10000000",
1659 => "10000000",
1660 => "10000000",
1661 => "10000000",
1662 => "10000000",
1663 => "10000000",
1664 => "10000000",
1665 => "10000000",
1666 => "10000000",
1667 => "10000000",
1668 => "10000000",
1669 => "10000000",
1670 => "10000000",
1671 => "10000000",
1672 => "10000000",
1673 => "10000000",
1674 => "10000000",
1675 => "10000000",
1676 => "10000000",
1677 => "10000000",
1678 => "10000000",
1679 => "10000000",
1680 => "10000000",
1681 => "10000000",
1682 => "10000000",
1683 => "10000000",
1684 => "10000000",
1685 => "10000000",
1686 => "10000000",
1687 => "10000000",
1688 => "10000000",
1689 => "10000000",
1690 => "10000000",
1691 => "10000000",
1692 => "10000000",
1693 => "10000000",
1694 => "10000000",
1695 => "10000000",
1696 => "10000000",
1697 => "10000000",
1698 => "10000000",
1699 => "10000000",
1700 => "10000000",
1701 => "10000000",
1702 => "10000000",
1703 => "10000000",
1704 => "10000000",
1705 => "10000000",
1706 => "10000000",
1707 => "10000000",
1708 => "10000000",
1709 => "10000000",
1710 => "10000000",
1711 => "10000000",
1712 => "10000000",
1713 => "10000000",
1714 => "10000000",
1715 => "10000000",
1716 => "10000000",
1717 => "10000000",
1718 => "10000000",
1719 => "10000000",
1720 => "11111111",
1721 => "00000001",
1722 => "00000001",
1723 => "11111111",
1724 => "10000000",
1725 => "10000000",
1726 => "10000000",
1727 => "10000000",
1728 => "10000000",
1729 => "10000000",
1730 => "10000000",
1731 => "10000000",
1732 => "10000000",
1733 => "10000000",
1734 => "10000000",
1735 => "10000000",
1736 => "10000000",
1737 => "10000000",
1738 => "10000000",
1739 => "10000000",
1740 => "10000000",
1741 => "10000000",
1742 => "10000000",
1743 => "10000000",
1744 => "10000000",
1745 => "10000000",
1746 => "10000000",
1747 => "10000000",
1748 => "10000000",
1749 => "10000000",
1750 => "10000000",
1751 => "10000000",
1752 => "10000000",
1753 => "10000000",
1754 => "10000000",
1755 => "10000000",
1756 => "10000000",
1757 => "10000000",
1758 => "10000000",
1759 => "10000000",
1760 => "10000000",
1761 => "10000000",
1762 => "10000000",
1763 => "10000000",
1764 => "10000000",
1765 => "10000000",
1766 => "10000000",
1767 => "10000000",
1768 => "10000000",
1769 => "10000000",
1770 => "10000000",
1771 => "10000000",
1772 => "10000000",
1773 => "10000000",
1774 => "10000000",
1775 => "10000000",
1776 => "10000000",
1777 => "10000000",
1778 => "10000000",
1779 => "10000000",
1780 => "10000000",
1781 => "10000000",
1782 => "10000000",
1783 => "10000000",
1784 => "10000000",
1785 => "10000000",
1786 => "10000000",
1787 => "10000000",
1788 => "10000000",
1789 => "10000000",
1790 => "10000000",
1791 => "10000000",
1792 => "10000000",
1793 => "10000000",
1794 => "10000000",
1795 => "10000000",
1796 => "10000000",
1797 => "10000000",
1798 => "10000000",
1799 => "10000000",
1800 => "10000000",
1801 => "10000000",
1802 => "11111111",
1803 => "00000001",
1804 => "00000001",
1805 => "11111111",
1806 => "10000000",
1807 => "10000000",
1808 => "10000000",
1809 => "10000000",
1810 => "10000000",
1811 => "10000000",
1812 => "10000000",
1813 => "10000000",
1814 => "10000000",
1815 => "10000000",
1816 => "10000000",
1817 => "10000000",
1818 => "10000000",
1819 => "10000000",
1820 => "10000000",
1821 => "10000000",
1822 => "10000000",
1823 => "10000000",
1824 => "10000000",
1825 => "10000000",
1826 => "10000000",
1827 => "10000000",
1828 => "10000000",
1829 => "10000000",
1830 => "10000000",
1831 => "10000000",
1832 => "10000000",
1833 => "10000000",
1834 => "10000000",
1835 => "10000000",
1836 => "10000000",
1837 => "10000000",
1838 => "10000000",
1839 => "10000000",
1840 => "10000000",
1841 => "10000000",
1842 => "10000000",
1843 => "10000000",
1844 => "10000000",
1845 => "10000000",
1846 => "10000000",
1847 => "10000000",
1848 => "10000000",
1849 => "10000000",
1850 => "10000000",
1851 => "10000000",
1852 => "10000000",
1853 => "10000000",
1854 => "10000000",
1855 => "10000000",
1856 => "10000000",
1857 => "10000000",
1858 => "10000000",
1859 => "10000000",
1860 => "10000000",
1861 => "10000000",
1862 => "10000000",
1863 => "10000000",
1864 => "10000000",
1865 => "10000000",
1866 => "10000000",
1867 => "10000000",
1868 => "10000000",
1869 => "10000000",
1870 => "10000000",
1871 => "10000000",
1872 => "10000000",
1873 => "10000000",
1874 => "10000000",
1875 => "10000000",
1876 => "10000000",
1877 => "10000000",
1878 => "10000000",
1879 => "10000000",
1880 => "10000000",
1881 => "10000000",
1882 => "10000000",
1883 => "10000000",
1884 => "11111111",
1885 => "00000001",
1886 => "00000001",
1887 => "11111111",
1888 => "10000000",
1889 => "10000000",
1890 => "10000000",
1891 => "10000000",
1892 => "10000000",
1893 => "10000000",
1894 => "10000000",
1895 => "10000000",
1896 => "10000000",
1897 => "10000000",
1898 => "10000000",
1899 => "10000000",
1900 => "10000000",
1901 => "10000000",
1902 => "10000000",
1903 => "10000000",
1904 => "10000000",
1905 => "10000000",
1906 => "10000000",
1907 => "10000000",
1908 => "10000000",
1909 => "10000000",
1910 => "10000000",
1911 => "10000000",
1912 => "10000000",
1913 => "10000000",
1914 => "10000000",
1915 => "10000000",
1916 => "10000000",
1917 => "10000000",
1918 => "10000000",
1919 => "10000000",
1920 => "10000000",
1921 => "10000000",
1922 => "10000000",
1923 => "10000000",
1924 => "10000000",
1925 => "10000000",
1926 => "10000000",
1927 => "10000000",
1928 => "10000000",
1929 => "10000000",
1930 => "10000000",
1931 => "10000000",
1932 => "10000000",
1933 => "10000000",
1934 => "10000000",
1935 => "10000000",
1936 => "10000000",
1937 => "10000000",
1938 => "10000000",
1939 => "10000000",
1940 => "10000000",
1941 => "10000000",
1942 => "10000000",
1943 => "10000000",
1944 => "10000000",
1945 => "10000000",
1946 => "10000000",
1947 => "10000000",
1948 => "10000000",
1949 => "10000000",
1950 => "10000000",
1951 => "10000000",
1952 => "10000000",
1953 => "10000000",
1954 => "10000000",
1955 => "10000000",
1956 => "10000000",
1957 => "10000000",
1958 => "10000000",
1959 => "10000000",
1960 => "10000000",
1961 => "10000000",
1962 => "10000000",
1963 => "10000000",
1964 => "10000000",
1965 => "10000000",
1966 => "11111111",
1967 => "00000001",
1968 => "00000001",
1969 => "11111111",
1970 => "10000000",
1971 => "10000000",
1972 => "10000000",
1973 => "10000000",
1974 => "10000000",
1975 => "10000000",
1976 => "10000000",
1977 => "10000000",
1978 => "10000000",
1979 => "10000000",
1980 => "10000000",
1981 => "10000000",
1982 => "10000000",
1983 => "10000000",
1984 => "10000000",
1985 => "10000000",
1986 => "10000000",
1987 => "10000000",
1988 => "10000000",
1989 => "10000000",
1990 => "10000000",
1991 => "10000000",
1992 => "10000000",
1993 => "10000000",
1994 => "10000000",
1995 => "10000000",
1996 => "10000000",
1997 => "10000000",
1998 => "10000000",
1999 => "10000000",
2000 => "10000000",
2001 => "10000000",
2002 => "10000000",
2003 => "10000000",
2004 => "10000000",
2005 => "10000000",
2006 => "10000000",
2007 => "10000000",
2008 => "10000000",
2009 => "10000000",
2010 => "10000000",
2011 => "10000000",
2012 => "10000000",
2013 => "10000000",
2014 => "10000000",
2015 => "10000000",
2016 => "10000000",
2017 => "10000000",
2018 => "10000000",
2019 => "10000000",
2020 => "10000000",
2021 => "10000000",
2022 => "10000000",
2023 => "10000000",
2024 => "10000000",
2025 => "10000000",
2026 => "10000000",
2027 => "10000000",
2028 => "10000000",
2029 => "10000000",
2030 => "10000000",
2031 => "10000000",
2032 => "10000000",
2033 => "10000000",
2034 => "10000000",
2035 => "10000000",
2036 => "10000000",
2037 => "10000000",
2038 => "10000000",
2039 => "10000000",
2040 => "10000000",
2041 => "10000000",
2042 => "10000000",
2043 => "10000000",
2044 => "10000000",
2045 => "10000000",
2046 => "10000000",
2047 => "10000000",
2048 => "11111111",
2049 => "00000001",
2050 => "00000001",
2051 => "11111111",
2052 => "10000000",
2053 => "10000000",
2054 => "10000000",
2055 => "10000000",
2056 => "10000000",
2057 => "10000000",
2058 => "10000000",
2059 => "10000000",
2060 => "10000000",
2061 => "10000000",
2062 => "10000000",
2063 => "10000000",
2064 => "10000000",
2065 => "10000000",
2066 => "10000000",
2067 => "10000000",
2068 => "10000000",
2069 => "10000000",
2070 => "10000000",
2071 => "10000000",
2072 => "10000000",
2073 => "10000000",
2074 => "10000000",
2075 => "10000000",
2076 => "10000000",
2077 => "10000000",
2078 => "10000000",
2079 => "10000000",
2080 => "10000000",
2081 => "10000000",
2082 => "10000000",
2083 => "10000000",
2084 => "10000000",
2085 => "10000000",
2086 => "10000000",
2087 => "10000000",
2088 => "10000000",
2089 => "10000000",
2090 => "10000000",
2091 => "10000000",
2092 => "10000000",
2093 => "10000000",
2094 => "10000000",
2095 => "10000000",
2096 => "10000000",
2097 => "10000000",
2098 => "10000000",
2099 => "10000000",
2100 => "10000000",
2101 => "10000000",
2102 => "10000000",
2103 => "10000000",
2104 => "10000000",
2105 => "10000000",
2106 => "10000000",
2107 => "10000000",
2108 => "10000000",
2109 => "10000000",
2110 => "10000000",
2111 => "10000000",
2112 => "10000000",
2113 => "10000000",
2114 => "10000000",
2115 => "10000000",
2116 => "10000000",
2117 => "10000000",
2118 => "10000000",
2119 => "10000000",
2120 => "10000000",
2121 => "10000000",
2122 => "10000000",
2123 => "10000000",
2124 => "10000000",
2125 => "10000000",
2126 => "10000000",
2127 => "10000000",
2128 => "10000000",
2129 => "10000000",
2130 => "11111111",
2131 => "00000001",
2132 => "00000001",
2133 => "11111111",
2134 => "10000000",
2135 => "10000000",
2136 => "10000000",
2137 => "10000000",
2138 => "10000000",
2139 => "10000000",
2140 => "10000000",
2141 => "10000000",
2142 => "10000000",
2143 => "10000000",
2144 => "10000000",
2145 => "10000000",
2146 => "10000000",
2147 => "10000000",
2148 => "10000000",
2149 => "10000000",
2150 => "10000000",
2151 => "10000000",
2152 => "10000000",
2153 => "10000000",
2154 => "10000000",
2155 => "10000000",
2156 => "10000000",
2157 => "10000000",
2158 => "10000000",
2159 => "10000000",
2160 => "10000000",
2161 => "10000000",
2162 => "10000000",
2163 => "10000000",
2164 => "10000000",
2165 => "10000000",
2166 => "10000000",
2167 => "10000000",
2168 => "10000000",
2169 => "10000000",
2170 => "10000000",
2171 => "10000000",
2172 => "10000000",
2173 => "10000000",
2174 => "10000000",
2175 => "10000000",
2176 => "10000000",
2177 => "10000000",
2178 => "10000000",
2179 => "10000000",
2180 => "10000000",
2181 => "10000000",
2182 => "10000000",
2183 => "10000000",
2184 => "10000000",
2185 => "10000000",
2186 => "10000000",
2187 => "10000000",
2188 => "10000000",
2189 => "10000000",
2190 => "10000000",
2191 => "10000000",
2192 => "10000000",
2193 => "10000000",
2194 => "10000000",
2195 => "10000000",
2196 => "10000000",
2197 => "10000000",
2198 => "10000000",
2199 => "10000000",
2200 => "10000000",
2201 => "10000000",
2202 => "10000000",
2203 => "10000000",
2204 => "10000000",
2205 => "10000000",
2206 => "10000000",
2207 => "10000000",
2208 => "10000000",
2209 => "10000000",
2210 => "10000000",
2211 => "10000000",
2212 => "11111111",
2213 => "00000001",
2214 => "00000001",
2215 => "11111111",
2216 => "10000000",
2217 => "10000000",
2218 => "10000000",
2219 => "10000000",
2220 => "10000000",
2221 => "10000000",
2222 => "10000000",
2223 => "10000000",
2224 => "10000000",
2225 => "10000000",
2226 => "10000000",
2227 => "10000000",
2228 => "10000000",
2229 => "10000000",
2230 => "10000000",
2231 => "10000000",
2232 => "10000000",
2233 => "10000000",
2234 => "10000000",
2235 => "10000000",
2236 => "10000000",
2237 => "10000000",
2238 => "10000000",
2239 => "10000000",
2240 => "10000000",
2241 => "10000000",
2242 => "10000000",
2243 => "10000000",
2244 => "10000000",
2245 => "10000000",
2246 => "10000000",
2247 => "10000000",
2248 => "10000000",
2249 => "10000000",
2250 => "10000000",
2251 => "10000000",
2252 => "10000000",
2253 => "10000000",
2254 => "10000000",
2255 => "10000000",
2256 => "10000000",
2257 => "10000000",
2258 => "10000000",
2259 => "10000000",
2260 => "10000000",
2261 => "10000000",
2262 => "10000000",
2263 => "10000000",
2264 => "10000000",
2265 => "10000000",
2266 => "10000000",
2267 => "10000000",
2268 => "10000000",
2269 => "10000000",
2270 => "10000000",
2271 => "10000000",
2272 => "10000000",
2273 => "10000000",
2274 => "10000000",
2275 => "10000000",
2276 => "10000000",
2277 => "10000000",
2278 => "10000000",
2279 => "10000000",
2280 => "10000000",
2281 => "10000000",
2282 => "10000000",
2283 => "10000000",
2284 => "10000000",
2285 => "10000000",
2286 => "10000000",
2287 => "10000000",
2288 => "10000000",
2289 => "10000000",
2290 => "10000000",
2291 => "10000000",
2292 => "10000000",
2293 => "10000000",
2294 => "11111111",
2295 => "00000001",
2296 => "00000001",
2297 => "10110110",
2298 => "10101001",
2299 => "10000000",
2300 => "10000000",
2301 => "10000000",
2302 => "10000000",
2303 => "10000000",
2304 => "10000000",
2305 => "10000000",
2306 => "10000000",
2307 => "10000000",
2308 => "10000000",
2309 => "10000000",
2310 => "10000000",
2311 => "10000000",
2312 => "10000000",
2313 => "10000000",
2314 => "10000000",
2315 => "10000000",
2316 => "10000000",
2317 => "10000000",
2318 => "10000000",
2319 => "10000000",
2320 => "10000000",
2321 => "10000000",
2322 => "10000000",
2323 => "10000000",
2324 => "10000000",
2325 => "10000000",
2326 => "10000000",
2327 => "10000000",
2328 => "10000000",
2329 => "10000000",
2330 => "10000000",
2331 => "10000000",
2332 => "10000000",
2333 => "10000000",
2334 => "10000000",
2335 => "10000000",
2336 => "10000000",
2337 => "10000000",
2338 => "10000000",
2339 => "10000000",
2340 => "10000000",
2341 => "10000000",
2342 => "10000000",
2343 => "10000000",
2344 => "10000000",
2345 => "10000000",
2346 => "10000000",
2347 => "10000000",
2348 => "10000000",
2349 => "10000000",
2350 => "10000000",
2351 => "10000000",
2352 => "10000000",
2353 => "10000000",
2354 => "10000000",
2355 => "10000000",
2356 => "10000000",
2357 => "10000000",
2358 => "10000000",
2359 => "10000000",
2360 => "10000000",
2361 => "10000000",
2362 => "10000000",
2363 => "10000000",
2364 => "10000000",
2365 => "10000000",
2366 => "10000000",
2367 => "10000000",
2368 => "10000000",
2369 => "10000000",
2370 => "10000000",
2371 => "10000000",
2372 => "10000000",
2373 => "10000000",
2374 => "10000000",
2375 => "10101001",
2376 => "10110110",
2377 => "00000001",
2378 => "00000001",
2379 => "00100101",
2380 => "11111111",
2381 => "10101001",
2382 => "10000000",
2383 => "10000000",
2384 => "10000000",
2385 => "10000000",
2386 => "10000000",
2387 => "10000000",
2388 => "10000000",
2389 => "10000000",
2390 => "10000000",
2391 => "10000000",
2392 => "10000000",
2393 => "10000000",
2394 => "10000000",
2395 => "10000000",
2396 => "10000000",
2397 => "10000000",
2398 => "10000000",
2399 => "10000000",
2400 => "10000000",
2401 => "10000000",
2402 => "10000000",
2403 => "10000000",
2404 => "10000000",
2405 => "10000000",
2406 => "10000000",
2407 => "10000000",
2408 => "10000000",
2409 => "10000000",
2410 => "10000000",
2411 => "10000000",
2412 => "10000000",
2413 => "10000000",
2414 => "10000000",
2415 => "10000000",
2416 => "10000000",
2417 => "10000000",
2418 => "10000000",
2419 => "10000000",
2420 => "10000000",
2421 => "10000000",
2422 => "10000000",
2423 => "10000000",
2424 => "10000000",
2425 => "10000000",
2426 => "10000000",
2427 => "10000000",
2428 => "10000000",
2429 => "10000000",
2430 => "10000000",
2431 => "10000000",
2432 => "10000000",
2433 => "10000000",
2434 => "10000000",
2435 => "10000000",
2436 => "10000000",
2437 => "10000000",
2438 => "10000000",
2439 => "10000000",
2440 => "10000000",
2441 => "10000000",
2442 => "10000000",
2443 => "10000000",
2444 => "10000000",
2445 => "10000000",
2446 => "10000000",
2447 => "10000000",
2448 => "10000000",
2449 => "10000000",
2450 => "10000000",
2451 => "10000000",
2452 => "10000000",
2453 => "10000000",
2454 => "10000000",
2455 => "10000000",
2456 => "10101001",
2457 => "11111111",
2458 => "00100101",
2459 => "00000001",
2460 => "00000001",
2461 => "00000001",
2462 => "00100101",
2463 => "10110110",
2464 => "11111111",
2465 => "11111111",
2466 => "11111111",
2467 => "11111111",
2468 => "11111111",
2469 => "11111111",
2470 => "11111111",
2471 => "11111111",
2472 => "11111111",
2473 => "11111111",
2474 => "11111111",
2475 => "11111111",
2476 => "11111111",
2477 => "11111111",
2478 => "11111111",
2479 => "11111111",
2480 => "11111111",
2481 => "11111111",
2482 => "11111111",
2483 => "11111111",
2484 => "11111111",
2485 => "11111111",
2486 => "11111111",
2487 => "11111111",
2488 => "11111111",
2489 => "11111111",
2490 => "11111111",
2491 => "11111111",
2492 => "11111111",
2493 => "11111111",
2494 => "11111111",
2495 => "11111111",
2496 => "11111111",
2497 => "11111111",
2498 => "11111111",
2499 => "11111111",
2500 => "11111111",
2501 => "11111111",
2502 => "11111111",
2503 => "11111111",
2504 => "11111111",
2505 => "11111111",
2506 => "11111111",
2507 => "11111111",
2508 => "11111111",
2509 => "11111111",
2510 => "11111111",
2511 => "11111111",
2512 => "11111111",
2513 => "11111111",
2514 => "11111111",
2515 => "11111111",
2516 => "11111111",
2517 => "11111111",
2518 => "11111111",
2519 => "11111111",
2520 => "11111111",
2521 => "11111111",
2522 => "11111111",
2523 => "11111111",
2524 => "11111111",
2525 => "11111111",
2526 => "11111111",
2527 => "11111111",
2528 => "11111111",
2529 => "11111111",
2530 => "11111111",
2531 => "11111111",
2532 => "11111111",
2533 => "11111111",
2534 => "11111111",
2535 => "11111111",
2536 => "11111111",
2537 => "11111111",
2538 => "10110110",
2539 => "00100101",
2540 => "00000001",
2541 => "00000001",
2542 => "00000001",
2543 => "00000001",
2544 => "00000001",
2545 => "00000001",
2546 => "00000001",
2547 => "00000001",
2548 => "00000001",
2549 => "00000001",
2550 => "00000001",
2551 => "00000001",
2552 => "00000001",
2553 => "00000001",
2554 => "00000001",
2555 => "00000001",
2556 => "00000001",
2557 => "00000001",
2558 => "00000001",
2559 => "00000001",
2560 => "00000001",
2561 => "00000001",
2562 => "00000001",
2563 => "00000001",
2564 => "00000001",
2565 => "00000001",
2566 => "00000001",
2567 => "00000001",
2568 => "00000001",
2569 => "00000001",
2570 => "00000001",
2571 => "00000001",
2572 => "00000001",
2573 => "00000001",
2574 => "00000001",
2575 => "00000001",
2576 => "00000001",
2577 => "00000001",
2578 => "00000001",
2579 => "00000001",
2580 => "00000001",
2581 => "00000001",
2582 => "00000001",
2583 => "00000001",
2584 => "00000001",
2585 => "00000001",
2586 => "00000001",
2587 => "00000001",
2588 => "00000001",
2589 => "00000001",
2590 => "00000001",
2591 => "00000001",
2592 => "00000001",
2593 => "00000001",
2594 => "00000001",
2595 => "00000001",
2596 => "00000001",
2597 => "00000001",
2598 => "00000001",
2599 => "00000001",
2600 => "00000001",
2601 => "00000001",
2602 => "00000001",
2603 => "00000001",
2604 => "00000001",
2605 => "00000001",
2606 => "00000001",
2607 => "00000001",
2608 => "00000001",
2609 => "00000001",
2610 => "00000001",
2611 => "00000001",
2612 => "00000001",
2613 => "00000001",
2614 => "00000001",
2615 => "00000001",
2616 => "00000001",
2617 => "00000001",
2618 => "00000001",
2619 => "00000001",
2620 => "00000001",
2621 => "00000001",
2622 => "00000001",
2623 => "00000001");
       
begin

    process(clk)
    begin
    
        if rising_edge(clk) then
                dout <= red(to_integer(unsigned(addr)));
        end if;
    end process;

end Behavioral;


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity Button_OneSec is
    port(clk, rst: in std_logic;
         addr: in std_logic_vector(9 downto 0);
         dout: out std_logic_vector(7 downto 0));
end Button_OneSec;

architecture Behavioral of Button_OneSec is

    type mem is array (0 to 755) of std_logic_vector(7 downto 0);
    signal One: mem := (
        0 => "00000001",
        1 => "00000001",
        2 => "00000001",
        3 => "00100101",
        4 => "01001001",
        5 => "01001001",
        6 => "01001001",
        7 => "01001001",
        8 => "01001001",
        9 => "01001001",
        10 => "01001001",
        11 => "01001001",
        12 => "01001001",
        13 => "01001001",
        14 => "01001001",
        15 => "01001001",
        16 => "01001001",
        17 => "01001001",
        18 => "01001001",
        19 => "01001001",
        20 => "01001001",
        21 => "01001001",
        22 => "01001001",
        23 => "00100001",
        24 => "00000001",
        25 => "00000001",
        26 => "00000001",
        27 => "00000001",
        28 => "00100101",
        29 => "10010010",
        30 => "11011011",
        31 => "11011111",
        32 => "11011111",
        33 => "11011111",
        34 => "11011111",
        35 => "11011111",
        36 => "11011111",
        37 => "11011111",
        38 => "11011111",
        39 => "11011111",
        40 => "11011111",
        41 => "11111111",
        42 => "11111111",
        43 => "11011111",
        44 => "11011111",
        45 => "11111111",
        46 => "11111111",
        47 => "11011111",
        48 => "11011111",
        49 => "11011011",
        50 => "10010011",
        51 => "01001010",
        52 => "00000001",
        53 => "00000001",
        54 => "00000001",
        55 => "01110010",
        56 => "11011111",
        57 => "10111110",
        58 => "10011010",
        59 => "10011001",
        60 => "10011010",
        61 => "10011010",
        62 => "10011001",
        63 => "10011001",
        64 => "10011001",
        65 => "10011101",
        66 => "10011110",
        67 => "10011010",
        68 => "10011010",
        69 => "10011001",
        70 => "10011001",
        71 => "10011110",
        72 => "10011010",
        73 => "10011010",
        74 => "10011001",
        75 => "10011010",
        76 => "10111110",
        77 => "11011111",
        78 => "10010111",
        79 => "00100101",
        80 => "00000001",
        81 => "00101001",
        82 => "10111011",
        83 => "10111110",
        84 => "01010000",
        85 => "00010000",
        86 => "00010000",
        87 => "00010000",
        88 => "00010000",
        89 => "00010000",
        90 => "00010000",
        91 => "00010000",
        92 => "00010000",
        93 => "00010000",
        94 => "00010000",
        95 => "00010000",
        96 => "00010000",
        97 => "00010000",
        98 => "00010000",
        99 => "00001100",
        100 => "00010000",
        101 => "00010000",
        102 => "00010000",
        103 => "00110000",
        104 => "10011010",
        105 => "11011111",
        106 => "01101110",
        107 => "00000001",
        108 => "01001001",
        109 => "11011111",
        110 => "10011010",
        111 => "00010000",
        112 => "00010000",
        113 => "00010000",
        114 => "00010000",
        115 => "00010000",
        116 => "00010000",
        117 => "00010000",
        118 => "00010000",
        119 => "00010000",
        120 => "00010000",
        121 => "00010000",
        122 => "00010000",
        123 => "00010000",
        124 => "00010000",
        125 => "00010000",
        126 => "00010000",
        127 => "00010000",
        128 => "00010000",
        129 => "00010000",
        130 => "00010000",
        131 => "01110101",
        132 => "11011111",
        133 => "10010010",
        134 => "00000001",
        135 => "01001001",
        136 => "11011111",
        137 => "01111001",
        138 => "00010000",
        139 => "00010000",
        140 => "00010000",
        141 => "00010000",
        142 => "00010000",
        143 => "00010000",
        144 => "00010000",
        145 => "00010000",
        146 => "00010000",
        147 => "00010000",
        148 => "00010000",
        149 => "00010000",
        150 => "00010000",
        151 => "00010000",
        152 => "00010000",
        153 => "00010100",
        154 => "00010000",
        155 => "00010000",
        156 => "00010000",
        157 => "00010000",
        158 => "01010101",
        159 => "11011111",
        160 => "10010010",
        161 => "00000000",
        162 => "01001001",
        163 => "11011111",
        164 => "01111001",
        165 => "00010000",
        166 => "00010000",
        167 => "00010000",
        168 => "00010000",
        169 => "00010000",
        170 => "00010000",
        171 => "00010000",
        172 => "00010000",
        173 => "00010000",
        174 => "00010000",
        175 => "00010000",
        176 => "00010000",
        177 => "00010100",
        178 => "00010100",
        179 => "00010000",
        180 => "00010000",
        181 => "00010000",
        182 => "00010000",
        183 => "00010000",
        184 => "00010000",
        185 => "01010101",
        186 => "11011111",
        187 => "10010010",
        188 => "00000001",
        189 => "01001001",
        190 => "11011111",
        191 => "01111001",
        192 => "00010000",
        193 => "00010000",
        194 => "00010000",
        195 => "00010000",
        196 => "00010000",
        197 => "00010000",
        198 => "00010000",
        199 => "00010000",
        200 => "00010000",
        201 => "00010000",
        202 => "00010000",
        203 => "00010000",
        204 => "00010000",
        205 => "00010000",
        206 => "00010000",
        207 => "00010000",
        208 => "00010000",
        209 => "00010000",
        210 => "00010000",
        211 => "00010000",
        212 => "01010101",
        213 => "11011111",
        214 => "10010010",
        215 => "00000001",
        216 => "01001001",
        217 => "11011111",
        218 => "10011001",
        219 => "00010000",
        220 => "00010000",
        221 => "00010000",
        222 => "00010000",
        223 => "00010000",
        224 => "00010000",
        225 => "00010000",
        226 => "00010000",
        227 => "00010000",
        228 => "00010000",
        229 => "00010000",
        230 => "00010000",
        231 => "00010000",
        232 => "00010000",
        233 => "00010000",
        234 => "00010000",
        235 => "00010000",
        236 => "00010000",
        237 => "00010000",
        238 => "00010000",
        239 => "01010101",
        240 => "11011111",
        241 => "10010010",
        242 => "00000001",
        243 => "01101010",
        244 => "11011111",
        245 => "10011001",
        246 => "00010000",
        247 => "00010000",
        248 => "00010000",
        249 => "00010000",
        250 => "00010000",
        251 => "00110100",
        252 => "00110100",
        253 => "00110100",
        254 => "00010000",
        255 => "00010000",
        256 => "00010000",
        257 => "00010000",
        258 => "00010000",
        259 => "00010000",
        260 => "00010000",
        261 => "00010000",
        262 => "00010000",
        263 => "00010000",
        264 => "00010000",
        265 => "00010000",
        266 => "01010101",
        267 => "11011111",
        268 => "10010010",
        269 => "00000001",
        270 => "01001001",
        271 => "11011111",
        272 => "01111001",
        273 => "00010000",
        274 => "00010000",
        275 => "00010000",
        276 => "00010000",
        277 => "00010100",
        278 => "01111001",
        279 => "10111110",
        280 => "10011101",
        281 => "00110000",
        282 => "00010000",
        283 => "00010000",
        284 => "00010000",
        285 => "00010000",
        286 => "00010000",
        287 => "00010000",
        288 => "00010000",
        289 => "00010000",
        290 => "00010000",
        291 => "00010000",
        292 => "00010000",
        293 => "01010101",
        294 => "11011111",
        295 => "10010010",
        296 => "00000001",
        297 => "01001001",
        298 => "11011111",
        299 => "01111001",
        300 => "00010000",
        301 => "00010000",
        302 => "00010000",
        303 => "00010100",
        304 => "01011101",
        305 => "10111110",
        306 => "11011110",
        307 => "10111001",
        308 => "00110000",
        309 => "00010000",
        310 => "00010000",
        311 => "00010100",
        312 => "00110100",
        313 => "00110100",
        314 => "00110100",
        315 => "00010100",
        316 => "00010000",
        317 => "00010000",
        318 => "00010000",
        319 => "00010000",
        320 => "01010101",
        321 => "11011111",
        322 => "10010010",
        323 => "00000001",
        324 => "01001001",
        325 => "11011111",
        326 => "10011001",
        327 => "00010000",
        328 => "00010000",
        329 => "00010000",
        330 => "00010100",
        331 => "01011001",
        332 => "01111001",
        333 => "10111110",
        334 => "10011001",
        335 => "00110000",
        336 => "00010000",
        337 => "00010000",
        338 => "01111001",
        339 => "10111110",
        340 => "10011101",
        341 => "01111101",
        342 => "01010100",
        343 => "00010000",
        344 => "00010000",
        345 => "00010000",
        346 => "00010000",
        347 => "01010101",
        348 => "11011111",
        349 => "10010010",
        350 => "00000001",
        351 => "01001001",
        352 => "11011111",
        353 => "10011001",
        354 => "00010000",
        355 => "00010000",
        356 => "00010000",
        357 => "00010000",
        358 => "00010000",
        359 => "01010101",
        360 => "10111110",
        361 => "10011001",
        362 => "00110000",
        363 => "00010000",
        364 => "00110100",
        365 => "10011110",
        366 => "10111110",
        367 => "01110101",
        368 => "00110000",
        369 => "00010000",
        370 => "00010000",
        371 => "00010000",
        372 => "00010000",
        373 => "00010000",
        374 => "01010101",
        375 => "11011111",
        376 => "10010010",
        377 => "00000001",
        378 => "01001001",
        379 => "11011111",
        380 => "01111001",
        381 => "00010000",
        382 => "00010000",
        383 => "00010000",
        384 => "00010000",
        385 => "00010000",
        386 => "01010100",
        387 => "10111110",
        388 => "10011001",
        389 => "00110000",
        390 => "00010000",
        391 => "00010000",
        392 => "01111001",
        393 => "10011110",
        394 => "11011110",
        395 => "10011001",
        396 => "01010100",
        397 => "00010000",
        398 => "00010000",
        399 => "00010000",
        400 => "00010000",
        401 => "01010101",
        402 => "11011111",
        403 => "10010010",
        404 => "00000001",
        405 => "01001001",
        406 => "11011111",
        407 => "01111001",
        408 => "00010000",
        409 => "00010000",
        410 => "00010000",
        411 => "00010000",
        412 => "00010000",
        413 => "01010101",
        414 => "10111110",
        415 => "10011101",
        416 => "00110000",
        417 => "00010000",
        418 => "00010000",
        419 => "00010000",
        420 => "00110101",
        421 => "10011010",
        422 => "11011110",
        423 => "10011101",
        424 => "00110100",
        425 => "00010000",
        426 => "00010000",
        427 => "00010000",
        428 => "01010101",
        429 => "11011111",
        430 => "10010010",
        431 => "00000001",
        432 => "01001001",
        433 => "11011111",
        434 => "01111001",
        435 => "00010000",
        436 => "00010000",
        437 => "00010000",
        438 => "00010000",
        439 => "00110100",
        440 => "01111001",
        441 => "10111110",
        442 => "10111101",
        443 => "01110100",
        444 => "00110000",
        445 => "00010000",
        446 => "00110100",
        447 => "01010101",
        448 => "01111001",
        449 => "10111110",
        450 => "10011101",
        451 => "00110100",
        452 => "00010000",
        453 => "00010000",
        454 => "00010000",
        455 => "01010101",
        456 => "11011111",
        457 => "10010010",
        458 => "00000001",
        459 => "01001001",
        460 => "11011111",
        461 => "10011001",
        462 => "00010000",
        463 => "00010000",
        464 => "00010000",
        465 => "00010100",
        466 => "01011001",
        467 => "01111001",
        468 => "10011101",
        469 => "10011101",
        470 => "01111001",
        471 => "00110100",
        472 => "00110100",
        473 => "01011001",
        474 => "01111101",
        475 => "10011101",
        476 => "01111001",
        477 => "00110100",
        478 => "00010000",
        479 => "00010000",
        480 => "00010000",
        481 => "00010000",
        482 => "01010101",
        483 => "11011111",
        484 => "10010010",
        485 => "00000001",
        486 => "01001101",
        487 => "11011111",
        488 => "01111001",
        489 => "00010000",
        490 => "00010000",
        491 => "00010000",
        492 => "00010000",
        493 => "00010000",
        494 => "00010000",
        495 => "00010000",
        496 => "00010000",
        497 => "00010000",
        498 => "00010000",
        499 => "00010000",
        500 => "00010000",
        501 => "00010000",
        502 => "00010000",
        503 => "00010000",
        504 => "00010000",
        505 => "00010000",
        506 => "00010000",
        507 => "00010000",
        508 => "00010000",
        509 => "01011001",
        510 => "11011111",
        511 => "10010010",
        512 => "00000001",
        513 => "01001001",
        514 => "11011111",
        515 => "10011001",
        516 => "00010000",
        517 => "00010000",
        518 => "00010000",
        519 => "00010000",
        520 => "00010000",
        521 => "00010000",
        522 => "00010000",
        523 => "00010000",
        524 => "00010000",
        525 => "00010000",
        526 => "00010000",
        527 => "00010000",
        528 => "00010000",
        529 => "00010000",
        530 => "00010000",
        531 => "00010000",
        532 => "00010000",
        533 => "00010000",
        534 => "00010000",
        535 => "00010000",
        536 => "01010101",
        537 => "11011111",
        538 => "10010010",
        539 => "00000001",
        540 => "01001001",
        541 => "11011111",
        542 => "10011010",
        543 => "00010000",
        544 => "00010000",
        545 => "00010000",
        546 => "00010000",
        547 => "00010000",
        548 => "00010000",
        549 => "00010000",
        550 => "00010000",
        551 => "00010000",
        552 => "00010000",
        553 => "00010000",
        554 => "00010000",
        555 => "00010000",
        556 => "00010000",
        557 => "00010000",
        558 => "00010000",
        559 => "00010000",
        560 => "00010000",
        561 => "00010000",
        562 => "00010000",
        563 => "01010100",
        564 => "11011111",
        565 => "10010010",
        566 => "00000001",
        567 => "01001001",
        568 => "11011111",
        569 => "01111010",
        570 => "00010000",
        571 => "00010000",
        572 => "00010100",
        573 => "00010100",
        574 => "00010000",
        575 => "00010000",
        576 => "00010000",
        577 => "00010000",
        578 => "00010000",
        579 => "00010000",
        580 => "00010000",
        581 => "00010000",
        582 => "00010000",
        583 => "00010000",
        584 => "00010000",
        585 => "00010000",
        586 => "00010000",
        587 => "00010000",
        588 => "00010000",
        589 => "00010000",
        590 => "01010101",
        591 => "11011111",
        592 => "10010010",
        593 => "00000001",
        594 => "01001001",
        595 => "11011111",
        596 => "10011010",
        597 => "00010000",
        598 => "00010000",
        599 => "00010000",
        600 => "00010000",
        601 => "00010000",
        602 => "00010000",
        603 => "00010100",
        604 => "00010000",
        605 => "00010000",
        606 => "00010000",
        607 => "00010000",
        608 => "00010000",
        609 => "00010100",
        610 => "00010000",
        611 => "00010000",
        612 => "00010000",
        613 => "00010000",
        614 => "00010000",
        615 => "00010000",
        616 => "00010000",
        617 => "01110101",
        618 => "11011111",
        619 => "10010010",
        620 => "00000001",
        621 => "01001001",
        622 => "11011111",
        623 => "10011010",
        624 => "00110000",
        625 => "00010000",
        626 => "00010000",
        627 => "00010000",
        628 => "00010000",
        629 => "00010000",
        630 => "00010000",
        631 => "00010000",
        632 => "00010000",
        633 => "00010000",
        634 => "00010000",
        635 => "00010000",
        636 => "00010000",
        637 => "00010000",
        638 => "00010000",
        639 => "00010000",
        640 => "00010000",
        641 => "00010000",
        642 => "00010000",
        643 => "00110000",
        644 => "10011001",
        645 => "11011111",
        646 => "10001110",
        647 => "00000001",
        648 => "00100101",
        649 => "10110111",
        650 => "11011111",
        651 => "10011010",
        652 => "01010101",
        653 => "01010101",
        654 => "01010101",
        655 => "01010101",
        656 => "01010101",
        657 => "01010101",
        658 => "01010101",
        659 => "01010101",
        660 => "01010101",
        661 => "01010101",
        662 => "01010101",
        663 => "01010101",
        664 => "01010101",
        665 => "01010101",
        666 => "01010101",
        667 => "01010101",
        668 => "01010101",
        669 => "01010101",
        670 => "10011001",
        671 => "10111111",
        672 => "10111011",
        673 => "01000101",
        674 => "00000001",
        675 => "00000001",
        676 => "01001010",
        677 => "10110111",
        678 => "11011111",
        679 => "11011111",
        680 => "11011111",
        681 => "11011111",
        682 => "11011111",
        683 => "11011111",
        684 => "11011111",
        685 => "11011111",
        686 => "11011111",
        687 => "11011111",
        688 => "11011111",
        689 => "11011111",
        690 => "11011111",
        691 => "11011111",
        692 => "11011111",
        693 => "11011111",
        694 => "11011111",
        695 => "11011111",
        696 => "11011111",
        697 => "11011111",
        698 => "10111011",
        699 => "01101110",
        700 => "00000001",
        701 => "00000001",
        702 => "00000001",
        703 => "00000001",
        704 => "00100110",
        705 => "01101110",
        706 => "10010010",
        707 => "10010010",
        708 => "10010010",
        709 => "10010010",
        710 => "10010010",
        711 => "10010010",
        712 => "10010011",
        713 => "10010011",
        714 => "10010011",
        715 => "10010011",
        716 => "10010010",
        717 => "10010010",
        718 => "10010010",
        719 => "10010010",
        720 => "10010110",
        721 => "10010010",
        722 => "10010010",
        723 => "10010110",
        724 => "01110010",
        725 => "01001010",
        726 => "00000001",
        727 => "00000001",
        728 => "00000001",
        729 => "00000001",
        730 => "00000001",
        731 => "00000001",
        732 => "00000001",
        733 => "00000001",
        734 => "00000000",
        735 => "00000000",
        736 => "00000000",
        737 => "00000000",
        738 => "00000000",
        739 => "00000000",
        740 => "00000001",
        741 => "00000001",
        742 => "00000000",
        743 => "00000000",
        744 => "00000000",
        745 => "00000000",
        746 => "00000000",
        747 => "00000000",
        748 => "00000000",
        749 => "00000000",
        750 => "00000000",
        751 => "00000001",
        752 => "00000001",
        753 => "00000001",
        754 => "00000001",
        755 => "00000001");
        
begin

    process(clk)
    begin
    
        if rising_edge(clk) then
            if rst = '1' then
                One <= (others => (others => '0'));
            else
                dout <= One(to_integer(unsigned(addr)));
            end if;
        end if;
    end process;

end Behavioral;

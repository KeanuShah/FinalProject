

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity YellowClass is
    port(clk: in std_logic;
         addr: in std_logic_vector(11 downto 0);
         dout: out std_logic_vector(7 downto 0));
end YellowClass;

architecture Behavioral of YellowClass is

    type mem is array (0 to 2623) of std_logic_vector(7 downto 0);
    signal Yellow: mem := (
            0 => "00000001",
1 => "00000001",
2 => "00000001",
3 => "00000001",
4 => "00000001",
5 => "00000001",
6 => "00000001",
7 => "00000001",
8 => "00000001",
9 => "00000001",
10 => "00000001",
11 => "00000001",
12 => "00000001",
13 => "00000001",
14 => "00000001",
15 => "00000001",
16 => "00000001",
17 => "00000001",
18 => "00000001",
19 => "00000001",
20 => "00000001",
21 => "00000001",
22 => "00000001",
23 => "00000001",
24 => "00000001",
25 => "00000001",
26 => "00000001",
27 => "00000001",
28 => "00000001",
29 => "00000001",
30 => "00000001",
31 => "00000001",
32 => "00000001",
33 => "00000001",
34 => "00000001",
35 => "00000001",
36 => "00000001",
37 => "00000001",
38 => "00000001",
39 => "00000001",
40 => "00000001",
41 => "00000001",
42 => "00000001",
43 => "00000001",
44 => "00000001",
45 => "00000001",
46 => "00000001",
47 => "00000001",
48 => "00000001",
49 => "00000001",
50 => "00000001",
51 => "00000001",
52 => "00000001",
53 => "00000001",
54 => "00000001",
55 => "00000001",
56 => "00000001",
57 => "00000001",
58 => "00000001",
59 => "00000001",
60 => "00000001",
61 => "00000001",
62 => "00000001",
63 => "00000001",
64 => "00000001",
65 => "00000001",
66 => "00000001",
67 => "00000001",
68 => "00000001",
69 => "00000001",
70 => "00000001",
71 => "00000001",
72 => "00000001",
73 => "00000001",
74 => "00000001",
75 => "00000001",
76 => "00000001",
77 => "00000001",
78 => "00000001",
79 => "00000001",
80 => "00000001",
81 => "00000001",
82 => "00000001",
83 => "00000001",
84 => "00100101",
85 => "10110110",
86 => "11111111",
87 => "11111111",
88 => "11111111",
89 => "11111111",
90 => "11111111",
91 => "11111111",
92 => "11111111",
93 => "11111111",
94 => "11111111",
95 => "11111111",
96 => "11111111",
97 => "11111111",
98 => "11111111",
99 => "11111111",
100 => "11111111",
101 => "11111111",
102 => "11111111",
103 => "11111111",
104 => "11111111",
105 => "11111111",
106 => "11111111",
107 => "11111111",
108 => "11111111",
109 => "11111111",
110 => "11111111",
111 => "11111111",
112 => "11111111",
113 => "11111111",
114 => "11111111",
115 => "11111111",
116 => "11111111",
117 => "11111111",
118 => "11111111",
119 => "11111111",
120 => "11111111",
121 => "11111111",
122 => "11111111",
123 => "11111111",
124 => "11111111",
125 => "11111111",
126 => "11111111",
127 => "11111111",
128 => "11111111",
129 => "11111111",
130 => "11111111",
131 => "11111111",
132 => "11111111",
133 => "11111111",
134 => "11111111",
135 => "11111111",
136 => "11111111",
137 => "11111111",
138 => "11111111",
139 => "11111111",
140 => "11111111",
141 => "11111111",
142 => "11111111",
143 => "11111111",
144 => "11111111",
145 => "11111111",
146 => "11111111",
147 => "11111111",
148 => "11111111",
149 => "11111111",
150 => "11111111",
151 => "11111111",
152 => "11111111",
153 => "11111111",
154 => "11111111",
155 => "11111111",
156 => "11111111",
157 => "11111111",
158 => "11111111",
159 => "11111111",
160 => "10110110",
161 => "00100101",
162 => "00000001",
163 => "00000001",
164 => "00000001",
165 => "00100101",
166 => "11111111",
167 => "10110101",
168 => "10010000",
169 => "10010000",
170 => "10010000",
171 => "10010000",
172 => "10010000",
173 => "10010000",
174 => "10010000",
175 => "10010000",
176 => "10010000",
177 => "10010000",
178 => "10010000",
179 => "10010000",
180 => "10010000",
181 => "10010000",
182 => "10010000",
183 => "10010000",
184 => "10010000",
185 => "10010000",
186 => "10010000",
187 => "10010000",
188 => "10010000",
189 => "10010000",
190 => "10010000",
191 => "10010000",
192 => "10010000",
193 => "10010000",
194 => "10010000",
195 => "10010000",
196 => "10010000",
197 => "10010000",
198 => "10010000",
199 => "10010000",
200 => "10010000",
201 => "10010000",
202 => "10010000",
203 => "10010000",
204 => "10010000",
205 => "10010000",
206 => "10010000",
207 => "10010000",
208 => "10010000",
209 => "10010000",
210 => "10010000",
211 => "10010000",
212 => "10010000",
213 => "10010000",
214 => "10010000",
215 => "10010000",
216 => "10010000",
217 => "10010000",
218 => "10010000",
219 => "10010000",
220 => "10010000",
221 => "10010000",
222 => "10010000",
223 => "10010000",
224 => "10010000",
225 => "10010000",
226 => "10010000",
227 => "10010000",
228 => "10010000",
229 => "10010000",
230 => "10010000",
231 => "10010000",
232 => "10010000",
233 => "10010000",
234 => "10010000",
235 => "10010000",
236 => "10010000",
237 => "10010000",
238 => "10010000",
239 => "10010000",
240 => "10010000",
241 => "10010000",
242 => "10110101",
243 => "11111111",
244 => "00100101",
245 => "00000001",
246 => "00000001",
247 => "10110110",
248 => "10110101",
249 => "10010000",
250 => "10010000",
251 => "10010000",
252 => "10010000",
253 => "10010000",
254 => "10010000",
255 => "10010000",
256 => "10010000",
257 => "10010000",
258 => "10010000",
259 => "10010000",
260 => "10010000",
261 => "10010000",
262 => "10010000",
263 => "10010000",
264 => "10010000",
265 => "10010000",
266 => "10010000",
267 => "10010000",
268 => "10010000",
269 => "10010000",
270 => "10010000",
271 => "10010000",
272 => "10010000",
273 => "10010000",
274 => "10010000",
275 => "10010000",
276 => "10010000",
277 => "10010000",
278 => "10010000",
279 => "10010000",
280 => "10010000",
281 => "10010000",
282 => "10010000",
283 => "10010000",
284 => "10010000",
285 => "10010000",
286 => "10010000",
287 => "10010000",
288 => "10010000",
289 => "10010000",
290 => "10010000",
291 => "10010000",
292 => "10010000",
293 => "10010000",
294 => "10010000",
295 => "10010000",
296 => "10010000",
297 => "10010000",
298 => "10010000",
299 => "10010000",
300 => "10010000",
301 => "10010000",
302 => "10010000",
303 => "10010000",
304 => "10010000",
305 => "10010000",
306 => "10010000",
307 => "10010000",
308 => "10010000",
309 => "10010000",
310 => "10010000",
311 => "10010000",
312 => "10010000",
313 => "10010000",
314 => "10010000",
315 => "10010000",
316 => "10010000",
317 => "10010000",
318 => "10010000",
319 => "10010000",
320 => "10010000",
321 => "10010000",
322 => "10010000",
323 => "10010000",
324 => "10010000",
325 => "10110101",
326 => "10110110",
327 => "00000001",
328 => "00000001",
329 => "11111111",
330 => "10010000",
331 => "10010000",
332 => "10010000",
333 => "10010000",
334 => "10010000",
335 => "10010000",
336 => "10010000",
337 => "10010000",
338 => "10010000",
339 => "10010000",
340 => "10010000",
341 => "10010000",
342 => "10010000",
343 => "10010000",
344 => "10010000",
345 => "10010000",
346 => "10010000",
347 => "10010000",
348 => "10010000",
349 => "10010000",
350 => "10010000",
351 => "10010000",
352 => "10010000",
353 => "10010000",
354 => "10010000",
355 => "10010000",
356 => "10010000",
357 => "10010000",
358 => "10010000",
359 => "10010000",
360 => "10010000",
361 => "10010000",
362 => "10010000",
363 => "10010000",
364 => "10010000",
365 => "10010000",
366 => "10010000",
367 => "10010000",
368 => "10010000",
369 => "10010000",
370 => "10010000",
371 => "10010000",
372 => "10010000",
373 => "10010000",
374 => "10010000",
375 => "10010000",
376 => "10010000",
377 => "10010000",
378 => "10010000",
379 => "10010000",
380 => "10010000",
381 => "10010000",
382 => "10010000",
383 => "10010000",
384 => "10010000",
385 => "10010000",
386 => "10010000",
387 => "10010000",
388 => "10010000",
389 => "10010000",
390 => "10010000",
391 => "10010000",
392 => "10010000",
393 => "10010000",
394 => "10010000",
395 => "10010000",
396 => "10010000",
397 => "10010000",
398 => "10010000",
399 => "10010000",
400 => "10010000",
401 => "10010000",
402 => "10010000",
403 => "10010000",
404 => "10010000",
405 => "10010000",
406 => "10010000",
407 => "10010000",
408 => "11111111",
409 => "00000001",
410 => "00000001",
411 => "11111111",
412 => "10010000",
413 => "10010000",
414 => "10010000",
415 => "10010000",
416 => "10010000",
417 => "10010000",
418 => "10010000",
419 => "10010000",
420 => "10010000",
421 => "10010000",
422 => "10010000",
423 => "10010000",
424 => "10010000",
425 => "10010000",
426 => "10010000",
427 => "10010000",
428 => "10010000",
429 => "10010000",
430 => "10010000",
431 => "10010000",
432 => "10010000",
433 => "10010000",
434 => "10010000",
435 => "10010000",
436 => "10010000",
437 => "10010000",
438 => "10010000",
439 => "10010000",
440 => "10010000",
441 => "10010000",
442 => "10010000",
443 => "10010000",
444 => "10010000",
445 => "10010000",
446 => "10010000",
447 => "10010000",
448 => "10010000",
449 => "10010000",
450 => "10010000",
451 => "10010000",
452 => "10010000",
453 => "10010000",
454 => "10010000",
455 => "10010000",
456 => "10010000",
457 => "10010000",
458 => "10010000",
459 => "10010000",
460 => "10010000",
461 => "10010000",
462 => "10010000",
463 => "10010000",
464 => "10010000",
465 => "10010000",
466 => "10010000",
467 => "10010000",
468 => "10010000",
469 => "10010000",
470 => "10010000",
471 => "10010000",
472 => "10010000",
473 => "10010000",
474 => "10010000",
475 => "10010000",
476 => "10010000",
477 => "10010000",
478 => "10010000",
479 => "10010000",
480 => "10010000",
481 => "10010000",
482 => "10010000",
483 => "10010000",
484 => "10010000",
485 => "10010000",
486 => "10010000",
487 => "10010000",
488 => "10010000",
489 => "10010000",
490 => "11111111",
491 => "00000001",
492 => "00000001",
493 => "11111111",
494 => "10010000",
495 => "10010000",
496 => "10010000",
497 => "10010000",
498 => "10010000",
499 => "10010000",
500 => "10010000",
501 => "10010000",
502 => "10010000",
503 => "10010000",
504 => "10010000",
505 => "10010000",
506 => "10010000",
507 => "10010000",
508 => "10010000",
509 => "10010000",
510 => "10010000",
511 => "10010000",
512 => "10010000",
513 => "10010000",
514 => "10010000",
515 => "10010000",
516 => "10010000",
517 => "10010000",
518 => "10010000",
519 => "10010000",
520 => "10010000",
521 => "10010000",
522 => "10010000",
523 => "10010000",
524 => "10010000",
525 => "10010000",
526 => "10010000",
527 => "10010000",
528 => "10010000",
529 => "10010000",
530 => "10010000",
531 => "10010000",
532 => "10010000",
533 => "10010000",
534 => "10010000",
535 => "10010000",
536 => "10010000",
537 => "10010000",
538 => "10010000",
539 => "10010000",
540 => "10010000",
541 => "10010000",
542 => "10010000",
543 => "10010000",
544 => "10010000",
545 => "10010000",
546 => "10010000",
547 => "10010000",
548 => "10010000",
549 => "10010000",
550 => "10010000",
551 => "10010000",
552 => "10010000",
553 => "10010000",
554 => "10010000",
555 => "10010000",
556 => "10010000",
557 => "10010000",
558 => "10010000",
559 => "10010000",
560 => "10010000",
561 => "10010000",
562 => "10010000",
563 => "10010000",
564 => "10010000",
565 => "10010000",
566 => "10010000",
567 => "10010000",
568 => "10010000",
569 => "10010000",
570 => "10010000",
571 => "10010000",
572 => "11111111",
573 => "00000001",
574 => "00000001",
575 => "11111111",
576 => "10010000",
577 => "10010000",
578 => "10010000",
579 => "10010000",
580 => "10010000",
581 => "10010000",
582 => "10010000",
583 => "10010000",
584 => "10010000",
585 => "10010000",
586 => "10010000",
587 => "10010000",
588 => "10010000",
589 => "10010000",
590 => "10010000",
591 => "10010000",
592 => "10010000",
593 => "10010000",
594 => "10010000",
595 => "10010000",
596 => "10010000",
597 => "10010000",
598 => "10010000",
599 => "10010000",
600 => "10010000",
601 => "10010000",
602 => "10010000",
603 => "10010000",
604 => "10010000",
605 => "10010000",
606 => "10010000",
607 => "10010000",
608 => "10010000",
609 => "10010000",
610 => "10010000",
611 => "10010000",
612 => "10010000",
613 => "10010000",
614 => "10010000",
615 => "10010000",
616 => "10010000",
617 => "10010000",
618 => "10010000",
619 => "10010000",
620 => "10010000",
621 => "10010000",
622 => "10010000",
623 => "10010000",
624 => "10010000",
625 => "10010000",
626 => "10010000",
627 => "10010000",
628 => "10010000",
629 => "10010000",
630 => "10010000",
631 => "10010000",
632 => "10010000",
633 => "10010000",
634 => "10010000",
635 => "10010000",
636 => "10010000",
637 => "10010000",
638 => "10010000",
639 => "10010000",
640 => "10010000",
641 => "10010000",
642 => "10010000",
643 => "10010000",
644 => "10010000",
645 => "10010000",
646 => "10010000",
647 => "10010000",
648 => "10010000",
649 => "10010000",
650 => "10010000",
651 => "10010000",
652 => "10010000",
653 => "10010000",
654 => "11111111",
655 => "00000001",
656 => "00000001",
657 => "11111111",
658 => "10010000",
659 => "10010000",
660 => "10010000",
661 => "10010000",
662 => "10010000",
663 => "10010000",
664 => "10010000",
665 => "10010000",
666 => "10010000",
667 => "10010000",
668 => "10010000",
669 => "10010000",
670 => "10010000",
671 => "10010000",
672 => "10010000",
673 => "10010000",
674 => "10010000",
675 => "10010000",
676 => "10010000",
677 => "10010000",
678 => "10010000",
679 => "10010000",
680 => "10010000",
681 => "10010000",
682 => "10010000",
683 => "10010000",
684 => "10010000",
685 => "10010000",
686 => "10010000",
687 => "10010000",
688 => "10010000",
689 => "10010000",
690 => "10010000",
691 => "10010000",
692 => "10010000",
693 => "10010000",
694 => "10010000",
695 => "10010000",
696 => "10010000",
697 => "10010000",
698 => "10010000",
699 => "10010000",
700 => "10010000",
701 => "10010000",
702 => "10010000",
703 => "10010000",
704 => "10010000",
705 => "10010000",
706 => "10010000",
707 => "10010000",
708 => "10010000",
709 => "10010000",
710 => "10010000",
711 => "10010000",
712 => "10010000",
713 => "10010000",
714 => "10010000",
715 => "10010000",
716 => "10010000",
717 => "10010000",
718 => "10010000",
719 => "10010000",
720 => "10010000",
721 => "10010000",
722 => "10010000",
723 => "10010000",
724 => "10010000",
725 => "10010000",
726 => "10010000",
727 => "10010000",
728 => "10010000",
729 => "10010000",
730 => "10010000",
731 => "10010000",
732 => "10010000",
733 => "10010000",
734 => "10010000",
735 => "10010000",
736 => "11111111",
737 => "00000001",
738 => "00000001",
739 => "11111111",
740 => "10010000",
741 => "10010000",
742 => "10010000",
743 => "10010000",
744 => "10010000",
745 => "10010000",
746 => "10010000",
747 => "10010000",
748 => "10010000",
749 => "10010000",
750 => "10010000",
751 => "10010000",
752 => "10010000",
753 => "10010000",
754 => "10010000",
755 => "10010000",
756 => "10010000",
757 => "10010000",
758 => "10010000",
759 => "10010000",
760 => "10010000",
761 => "10010000",
762 => "10010000",
763 => "10010000",
764 => "10010000",
765 => "10010000",
766 => "10010000",
767 => "10010000",
768 => "10010000",
769 => "10010000",
770 => "10010000",
771 => "10010000",
772 => "10010000",
773 => "10010000",
774 => "10010000",
775 => "10010000",
776 => "10010000",
777 => "10010000",
778 => "10010000",
779 => "10010000",
780 => "10010000",
781 => "10010000",
782 => "10010000",
783 => "10010000",
784 => "10010000",
785 => "10010000",
786 => "10010000",
787 => "10010000",
788 => "10010000",
789 => "10010000",
790 => "10010000",
791 => "10010000",
792 => "10010000",
793 => "10010000",
794 => "10010000",
795 => "10010000",
796 => "10010000",
797 => "10010000",
798 => "10010000",
799 => "10010000",
800 => "10010000",
801 => "10010000",
802 => "10010000",
803 => "10010000",
804 => "10010000",
805 => "10010000",
806 => "10010000",
807 => "10010000",
808 => "10010000",
809 => "10010000",
810 => "10010000",
811 => "10010000",
812 => "10010000",
813 => "10010000",
814 => "10010000",
815 => "10010000",
816 => "10010000",
817 => "10010000",
818 => "11111111",
819 => "00000001",
820 => "00000001",
821 => "11111111",
822 => "10010000",
823 => "10010000",
824 => "10010000",
825 => "10010000",
826 => "10010000",
827 => "10010000",
828 => "10010000",
829 => "10010000",
830 => "10010000",
831 => "10010000",
832 => "10010000",
833 => "10010000",
834 => "10010000",
835 => "10010000",
836 => "10010000",
837 => "10010000",
838 => "10010000",
839 => "10010000",
840 => "10010000",
841 => "10010000",
842 => "10010000",
843 => "10010000",
844 => "10010000",
845 => "10010000",
846 => "10010000",
847 => "10010000",
848 => "10010000",
849 => "10010000",
850 => "10010000",
851 => "10010000",
852 => "10010000",
853 => "10010000",
854 => "10010000",
855 => "10010000",
856 => "10010000",
857 => "10010000",
858 => "10010000",
859 => "10010000",
860 => "10010000",
861 => "10010000",
862 => "10010000",
863 => "10010000",
864 => "10010000",
865 => "10010000",
866 => "10010000",
867 => "10010000",
868 => "10010000",
869 => "10010000",
870 => "10010000",
871 => "10010000",
872 => "10010000",
873 => "10010000",
874 => "10010000",
875 => "10010000",
876 => "10010000",
877 => "10010000",
878 => "10010000",
879 => "10010000",
880 => "10010000",
881 => "10010000",
882 => "10010000",
883 => "10010000",
884 => "10010000",
885 => "10010000",
886 => "10010000",
887 => "10010000",
888 => "10010000",
889 => "10010000",
890 => "10010000",
891 => "10010000",
892 => "10010000",
893 => "10010000",
894 => "10010000",
895 => "10010000",
896 => "10010000",
897 => "10010000",
898 => "10010000",
899 => "10010000",
900 => "11111111",
901 => "00000001",
902 => "00000001",
903 => "11111111",
904 => "10010000",
905 => "10010000",
906 => "10010000",
907 => "10010000",
908 => "10010000",
909 => "10010000",
910 => "10010000",
911 => "10010000",
912 => "10010000",
913 => "10010000",
914 => "10010000",
915 => "10010000",
916 => "10010000",
917 => "10010000",
918 => "10010000",
919 => "10010000",
920 => "10010000",
921 => "10010000",
922 => "10010000",
923 => "10010000",
924 => "10010000",
925 => "10010000",
926 => "10010000",
927 => "10010000",
928 => "10010000",
929 => "10010000",
930 => "10010000",
931 => "10010000",
932 => "10010000",
933 => "10010000",
934 => "10010000",
935 => "10010000",
936 => "10010000",
937 => "10010000",
938 => "10010000",
939 => "11011111",
940 => "11111111",
941 => "11011000",
942 => "10010000",
943 => "10010000",
944 => "10010000",
945 => "10010000",
946 => "10010000",
947 => "10010000",
948 => "10010000",
949 => "10010000",
950 => "10010000",
951 => "10010000",
952 => "10010000",
953 => "10010000",
954 => "10010000",
955 => "10010000",
956 => "10010000",
957 => "10010000",
958 => "10010000",
959 => "10010000",
960 => "10010000",
961 => "10010000",
962 => "10010000",
963 => "10010000",
964 => "10010000",
965 => "10010000",
966 => "10010000",
967 => "10010000",
968 => "10010000",
969 => "10010000",
970 => "10010000",
971 => "10010000",
972 => "10010000",
973 => "10010000",
974 => "10010000",
975 => "10010000",
976 => "10010000",
977 => "10010000",
978 => "10010000",
979 => "10010000",
980 => "10010000",
981 => "10010000",
982 => "11111111",
983 => "00000001",
984 => "00000001",
985 => "11111111",
986 => "10010000",
987 => "10010000",
988 => "10010000",
989 => "10010000",
990 => "10010000",
991 => "10010000",
992 => "10010000",
993 => "10010000",
994 => "10010000",
995 => "10010000",
996 => "10010000",
997 => "10010000",
998 => "10010000",
999 => "10010000",
1000 => "10010000",
1001 => "10010000",
1002 => "10010000",
1003 => "10010000",
1004 => "10010000",
1005 => "10010000",
1006 => "10010000",
1007 => "10010000",
1008 => "10010000",
1009 => "10010000",
1010 => "10010000",
1011 => "10010000",
1012 => "10010001",
1013 => "11111111",
1014 => "11111110",
1015 => "11010000",
1016 => "11011011",
1017 => "11111111",
1018 => "11111000",
1019 => "10010000",
1020 => "10010000",
1021 => "11011111",
1022 => "11111111",
1023 => "11011000",
1024 => "10010000",
1025 => "10010000",
1026 => "11011011",
1027 => "11111111",
1028 => "11111111",
1029 => "11111110",
1030 => "11010000",
1031 => "10010000",
1032 => "10010000",
1033 => "10010000",
1034 => "10010000",
1035 => "10010000",
1036 => "11011111",
1037 => "11111110",
1038 => "11010000",
1039 => "10010000",
1040 => "10010000",
1041 => "10010000",
1042 => "10010000",
1043 => "10010000",
1044 => "10010000",
1045 => "10010000",
1046 => "10010000",
1047 => "10010000",
1048 => "10010000",
1049 => "10010000",
1050 => "10010000",
1051 => "10010000",
1052 => "10010000",
1053 => "10010000",
1054 => "10010000",
1055 => "10010000",
1056 => "10010000",
1057 => "10010000",
1058 => "10010000",
1059 => "10010000",
1060 => "10010000",
1061 => "10010000",
1062 => "10010000",
1063 => "10010000",
1064 => "11111111",
1065 => "00000001",
1066 => "00000001",
1067 => "11111111",
1068 => "10010000",
1069 => "10010000",
1070 => "10010000",
1071 => "10010000",
1072 => "10010000",
1073 => "10010000",
1074 => "10010000",
1075 => "10010000",
1076 => "10010000",
1077 => "10010000",
1078 => "10010000",
1079 => "10010000",
1080 => "10010000",
1081 => "10010000",
1082 => "10010000",
1083 => "10010000",
1084 => "10010000",
1085 => "10010000",
1086 => "10010000",
1087 => "10010000",
1088 => "10010000",
1089 => "10010000",
1090 => "10010000",
1091 => "10010000",
1092 => "10010000",
1093 => "10010000",
1094 => "10010001",
1095 => "11111111",
1096 => "11111110",
1097 => "11010000",
1098 => "11011111",
1099 => "11111111",
1100 => "11111000",
1101 => "10010000",
1102 => "10010000",
1103 => "10010000",
1104 => "10010000",
1105 => "10010000",
1106 => "10010000",
1107 => "10010000",
1108 => "10010000",
1109 => "10010001",
1110 => "11011111",
1111 => "11111110",
1112 => "11010000",
1113 => "10010000",
1114 => "10010000",
1115 => "10010000",
1116 => "10010000",
1117 => "10010000",
1118 => "11011111",
1119 => "11111110",
1120 => "11010000",
1121 => "10010000",
1122 => "10010000",
1123 => "10010000",
1124 => "10010000",
1125 => "10010000",
1126 => "10010000",
1127 => "10010000",
1128 => "10010000",
1129 => "10010000",
1130 => "10010000",
1131 => "10010000",
1132 => "10010000",
1133 => "10010000",
1134 => "10010000",
1135 => "10010000",
1136 => "10010000",
1137 => "10010000",
1138 => "10010000",
1139 => "10010000",
1140 => "10010000",
1141 => "10010000",
1142 => "10010000",
1143 => "10010000",
1144 => "10010000",
1145 => "10010000",
1146 => "11111111",
1147 => "00000001",
1148 => "00000001",
1149 => "11111111",
1150 => "10010000",
1151 => "10010000",
1152 => "10010000",
1153 => "10010000",
1154 => "10010000",
1155 => "10010000",
1156 => "10010000",
1157 => "10010000",
1158 => "10010000",
1159 => "10010000",
1160 => "10010000",
1161 => "10010000",
1162 => "10010000",
1163 => "10010000",
1164 => "10010000",
1165 => "10010000",
1166 => "10010000",
1167 => "10010000",
1168 => "10010000",
1169 => "10010000",
1170 => "10010000",
1171 => "10010000",
1172 => "10010000",
1173 => "10010000",
1174 => "10010000",
1175 => "10010000",
1176 => "10011010",
1177 => "11111110",
1178 => "11111111",
1179 => "11011001",
1180 => "11111110",
1181 => "11111111",
1182 => "11111001",
1183 => "10011010",
1184 => "11111111",
1185 => "11111111",
1186 => "11111111",
1187 => "11011000",
1188 => "10010000",
1189 => "10010000",
1190 => "10010000",
1191 => "10010001",
1192 => "11011111",
1193 => "11111110",
1194 => "11010000",
1195 => "10010000",
1196 => "10010000",
1197 => "10011010",
1198 => "11111111",
1199 => "11111111",
1200 => "11111111",
1201 => "11111110",
1202 => "11010000",
1203 => "10010000",
1204 => "10010000",
1205 => "10010000",
1206 => "10010000",
1207 => "10010000",
1208 => "10010000",
1209 => "10010000",
1210 => "10010000",
1211 => "10010000",
1212 => "10010000",
1213 => "10010000",
1214 => "10010000",
1215 => "10010000",
1216 => "10010000",
1217 => "10010000",
1218 => "10010000",
1219 => "10010000",
1220 => "10010000",
1221 => "10010000",
1222 => "10010000",
1223 => "10010000",
1224 => "10010000",
1225 => "10010000",
1226 => "10010000",
1227 => "10010000",
1228 => "11111111",
1229 => "00000001",
1230 => "00000001",
1231 => "11111111",
1232 => "10010000",
1233 => "10010000",
1234 => "10010000",
1235 => "10010000",
1236 => "10010000",
1237 => "10010000",
1238 => "10010000",
1239 => "10010000",
1240 => "10010000",
1241 => "10010000",
1242 => "10010000",
1243 => "10010000",
1244 => "10010000",
1245 => "10010000",
1246 => "10010000",
1247 => "10010000",
1248 => "10010000",
1249 => "10010000",
1250 => "10010000",
1251 => "10010000",
1252 => "10010000",
1253 => "10010000",
1254 => "10010000",
1255 => "10010000",
1256 => "10010000",
1257 => "10010000",
1258 => "10011010",
1259 => "11111110",
1260 => "11011011",
1261 => "11111010",
1262 => "11111101",
1263 => "11011111",
1264 => "11111001",
1265 => "10010000",
1266 => "10010000",
1267 => "11011011",
1268 => "11111111",
1269 => "11011000",
1270 => "10010000",
1271 => "10010000",
1272 => "10010000",
1273 => "10010001",
1274 => "11011111",
1275 => "11111110",
1276 => "11010000",
1277 => "10010000",
1278 => "10011010",
1279 => "11111111",
1280 => "11111000",
1281 => "10010000",
1282 => "11011111",
1283 => "11111110",
1284 => "11010000",
1285 => "10010000",
1286 => "10010000",
1287 => "10010000",
1288 => "10010000",
1289 => "10010000",
1290 => "10010000",
1291 => "10010000",
1292 => "10010000",
1293 => "10010000",
1294 => "10010000",
1295 => "10010000",
1296 => "10010000",
1297 => "10010000",
1298 => "10010000",
1299 => "10010000",
1300 => "10010000",
1301 => "10010000",
1302 => "10010000",
1303 => "10010000",
1304 => "10010000",
1305 => "10010000",
1306 => "10010000",
1307 => "10010000",
1308 => "10010000",
1309 => "10010000",
1310 => "11111111",
1311 => "00000001",
1312 => "00000001",
1313 => "11111111",
1314 => "10010000",
1315 => "10010000",
1316 => "10010000",
1317 => "10010000",
1318 => "10010000",
1319 => "10010000",
1320 => "10010000",
1321 => "10010000",
1322 => "10010000",
1323 => "10010000",
1324 => "10010000",
1325 => "10010000",
1326 => "10010000",
1327 => "10010000",
1328 => "10010000",
1329 => "10010000",
1330 => "10010000",
1331 => "10010000",
1332 => "10010000",
1333 => "10010000",
1334 => "10010000",
1335 => "10010000",
1336 => "10010000",
1337 => "10010000",
1338 => "10010000",
1339 => "10010000",
1340 => "10011010",
1341 => "11111110",
1342 => "11011010",
1343 => "11111111",
1344 => "11111000",
1345 => "11011111",
1346 => "11111001",
1347 => "10010000",
1348 => "10010000",
1349 => "11011011",
1350 => "11111111",
1351 => "11011000",
1352 => "10010000",
1353 => "10010000",
1354 => "10010000",
1355 => "10010001",
1356 => "11011111",
1357 => "11111110",
1358 => "11010000",
1359 => "10010000",
1360 => "11011011",
1361 => "11111110",
1362 => "11010000",
1363 => "10010000",
1364 => "11011111",
1365 => "11111110",
1366 => "11010000",
1367 => "10010000",
1368 => "10010000",
1369 => "10010000",
1370 => "10010000",
1371 => "10010000",
1372 => "10010000",
1373 => "10010000",
1374 => "10010000",
1375 => "10010000",
1376 => "10010000",
1377 => "10010000",
1378 => "10010000",
1379 => "10010000",
1380 => "10010000",
1381 => "10010000",
1382 => "10010000",
1383 => "10010000",
1384 => "10010000",
1385 => "10010000",
1386 => "10010000",
1387 => "10010000",
1388 => "10010000",
1389 => "10010000",
1390 => "10010000",
1391 => "10010000",
1392 => "11111111",
1393 => "00000001",
1394 => "00000001",
1395 => "11111111",
1396 => "10010000",
1397 => "10010000",
1398 => "10010000",
1399 => "10010000",
1400 => "10010000",
1401 => "10010000",
1402 => "10010000",
1403 => "10010000",
1404 => "10010000",
1405 => "10010000",
1406 => "10010000",
1407 => "10010000",
1408 => "10010000",
1409 => "10010000",
1410 => "10010000",
1411 => "10010000",
1412 => "10010000",
1413 => "10010000",
1414 => "10010000",
1415 => "10010000",
1416 => "10010000",
1417 => "10010000",
1418 => "10010000",
1419 => "10010000",
1420 => "10010000",
1421 => "10010000",
1422 => "10011010",
1423 => "11111110",
1424 => "11010001",
1425 => "11111111",
1426 => "11011000",
1427 => "11011111",
1428 => "11111001",
1429 => "10010000",
1430 => "10010000",
1431 => "11011011",
1432 => "11111111",
1433 => "11011000",
1434 => "10010000",
1435 => "10010000",
1436 => "10010000",
1437 => "10010001",
1438 => "11011111",
1439 => "11111110",
1440 => "11010000",
1441 => "10010000",
1442 => "11011011",
1443 => "11111110",
1444 => "11010000",
1445 => "10010000",
1446 => "11011111",
1447 => "11111110",
1448 => "11010000",
1449 => "10010000",
1450 => "10010000",
1451 => "10010000",
1452 => "10010000",
1453 => "10010000",
1454 => "10010000",
1455 => "10010000",
1456 => "10010000",
1457 => "10010000",
1458 => "10010000",
1459 => "10010000",
1460 => "10010000",
1461 => "10010000",
1462 => "10010000",
1463 => "10010000",
1464 => "10010000",
1465 => "10010000",
1466 => "10010000",
1467 => "10010000",
1468 => "10010000",
1469 => "10010000",
1470 => "10010000",
1471 => "10010000",
1472 => "10010000",
1473 => "10010000",
1474 => "11111111",
1475 => "00000001",
1476 => "00000001",
1477 => "11111111",
1478 => "10010000",
1479 => "10010000",
1480 => "10010000",
1481 => "10010000",
1482 => "10010000",
1483 => "10010000",
1484 => "10010000",
1485 => "10010000",
1486 => "10010000",
1487 => "10010000",
1488 => "10010000",
1489 => "10010000",
1490 => "10010000",
1491 => "10010000",
1492 => "10010000",
1493 => "10010000",
1494 => "10010000",
1495 => "10010000",
1496 => "10010000",
1497 => "10010000",
1498 => "10010000",
1499 => "10010000",
1500 => "10010000",
1501 => "10010000",
1502 => "10010000",
1503 => "10010000",
1504 => "10011010",
1505 => "11111110",
1506 => "11010000",
1507 => "10010000",
1508 => "10010000",
1509 => "11011111",
1510 => "11111101",
1511 => "10010000",
1512 => "10010000",
1513 => "11011011",
1514 => "11111111",
1515 => "11011000",
1516 => "10010000",
1517 => "10010000",
1518 => "10010000",
1519 => "10010001",
1520 => "11011111",
1521 => "11111110",
1522 => "11010000",
1523 => "10010000",
1524 => "10011010",
1525 => "11111111",
1526 => "11011000",
1527 => "10011010",
1528 => "11111111",
1529 => "11111110",
1530 => "11010000",
1531 => "10010000",
1532 => "10010000",
1533 => "10010000",
1534 => "10010000",
1535 => "10010000",
1536 => "10010000",
1537 => "10010000",
1538 => "10010000",
1539 => "10010000",
1540 => "10010000",
1541 => "10010000",
1542 => "10010000",
1543 => "10010000",
1544 => "10010000",
1545 => "10010000",
1546 => "10010000",
1547 => "10010000",
1548 => "10010000",
1549 => "10010000",
1550 => "10010000",
1551 => "10010000",
1552 => "10010000",
1553 => "10010000",
1554 => "10010000",
1555 => "10010000",
1556 => "11111111",
1557 => "00000001",
1558 => "00000001",
1559 => "11111111",
1560 => "10010000",
1561 => "10010000",
1562 => "10010000",
1563 => "10010000",
1564 => "10010000",
1565 => "10010000",
1566 => "10010000",
1567 => "10010000",
1568 => "10010000",
1569 => "10010000",
1570 => "10010000",
1571 => "10010000",
1572 => "10010000",
1573 => "10010000",
1574 => "10010000",
1575 => "10010000",
1576 => "10010000",
1577 => "10010000",
1578 => "10010000",
1579 => "10010000",
1580 => "10010000",
1581 => "10010000",
1582 => "10010000",
1583 => "10010000",
1584 => "10010000",
1585 => "10010000",
1586 => "10011010",
1587 => "11111110",
1588 => "11010000",
1589 => "10010000",
1590 => "10010000",
1591 => "11011111",
1592 => "11111101",
1593 => "10011010",
1594 => "11111111",
1595 => "11111111",
1596 => "11111111",
1597 => "11111111",
1598 => "11111110",
1599 => "11010000",
1600 => "11011111",
1601 => "11111111",
1602 => "11111111",
1603 => "11111111",
1604 => "11111111",
1605 => "11111001",
1606 => "10010000",
1607 => "11011111",
1608 => "11111111",
1609 => "11111111",
1610 => "11111111",
1611 => "11111110",
1612 => "11010000",
1613 => "10010000",
1614 => "10010000",
1615 => "10010000",
1616 => "10010000",
1617 => "10010000",
1618 => "10010000",
1619 => "10010000",
1620 => "10010000",
1621 => "10010000",
1622 => "10010000",
1623 => "10010000",
1624 => "10010000",
1625 => "10010000",
1626 => "10010000",
1627 => "10010000",
1628 => "10010000",
1629 => "10010000",
1630 => "10010000",
1631 => "10010000",
1632 => "10010000",
1633 => "10010000",
1634 => "10010000",
1635 => "10010000",
1636 => "10010000",
1637 => "10010000",
1638 => "11111111",
1639 => "00000001",
1640 => "00000001",
1641 => "11111111",
1642 => "10010000",
1643 => "10010000",
1644 => "10010000",
1645 => "10010000",
1646 => "10010000",
1647 => "10010000",
1648 => "10010000",
1649 => "10010000",
1650 => "10010000",
1651 => "10010000",
1652 => "10010000",
1653 => "10010000",
1654 => "10010000",
1655 => "10010000",
1656 => "10010000",
1657 => "10010000",
1658 => "10010000",
1659 => "10010000",
1660 => "10010000",
1661 => "10010000",
1662 => "10010000",
1663 => "10010000",
1664 => "10010000",
1665 => "10010000",
1666 => "10010000",
1667 => "10010000",
1668 => "10010000",
1669 => "10010000",
1670 => "10010000",
1671 => "10010000",
1672 => "10010000",
1673 => "10010000",
1674 => "10010000",
1675 => "10010000",
1676 => "10010000",
1677 => "10010000",
1678 => "10010000",
1679 => "10010000",
1680 => "10010000",
1681 => "10010000",
1682 => "10010000",
1683 => "10010000",
1684 => "10010000",
1685 => "10010000",
1686 => "10010000",
1687 => "10010000",
1688 => "10010000",
1689 => "10010000",
1690 => "10010000",
1691 => "10010000",
1692 => "10010000",
1693 => "10010000",
1694 => "10010000",
1695 => "10010000",
1696 => "10010000",
1697 => "10010000",
1698 => "10010000",
1699 => "10010000",
1700 => "10010000",
1701 => "10010000",
1702 => "10010000",
1703 => "10010000",
1704 => "10010000",
1705 => "10010000",
1706 => "10010000",
1707 => "10010000",
1708 => "10010000",
1709 => "10010000",
1710 => "10010000",
1711 => "10010000",
1712 => "10010000",
1713 => "10010000",
1714 => "10010000",
1715 => "10010000",
1716 => "10010000",
1717 => "10010000",
1718 => "10010000",
1719 => "10010000",
1720 => "11111111",
1721 => "00000001",
1722 => "00000001",
1723 => "11111111",
1724 => "10010000",
1725 => "10010000",
1726 => "10010000",
1727 => "10010000",
1728 => "10010000",
1729 => "10010000",
1730 => "10010000",
1731 => "10010000",
1732 => "10010000",
1733 => "10010000",
1734 => "10010000",
1735 => "10010000",
1736 => "10010000",
1737 => "10010000",
1738 => "10010000",
1739 => "10010000",
1740 => "10010000",
1741 => "10010000",
1742 => "10010000",
1743 => "10010000",
1744 => "10010000",
1745 => "10010000",
1746 => "10010000",
1747 => "10010000",
1748 => "10010000",
1749 => "10010000",
1750 => "10010000",
1751 => "10010000",
1752 => "10010000",
1753 => "10010000",
1754 => "10010000",
1755 => "10010000",
1756 => "10010000",
1757 => "10010000",
1758 => "10010000",
1759 => "10010000",
1760 => "10010000",
1761 => "10010000",
1762 => "10010000",
1763 => "10010000",
1764 => "10010000",
1765 => "10010000",
1766 => "10010000",
1767 => "10010000",
1768 => "10010000",
1769 => "10010000",
1770 => "10010000",
1771 => "10010000",
1772 => "10010000",
1773 => "10010000",
1774 => "10010000",
1775 => "10010000",
1776 => "10010000",
1777 => "10010000",
1778 => "10010000",
1779 => "10010000",
1780 => "10010000",
1781 => "10010000",
1782 => "10010000",
1783 => "10010000",
1784 => "10010000",
1785 => "10010000",
1786 => "10010000",
1787 => "10010000",
1788 => "10010000",
1789 => "10010000",
1790 => "10010000",
1791 => "10010000",
1792 => "10010000",
1793 => "10010000",
1794 => "10010000",
1795 => "10010000",
1796 => "10010000",
1797 => "10010000",
1798 => "10010000",
1799 => "10010000",
1800 => "10010000",
1801 => "10010000",
1802 => "11111111",
1803 => "00000001",
1804 => "00000001",
1805 => "11111111",
1806 => "10010000",
1807 => "10010000",
1808 => "10010000",
1809 => "10010000",
1810 => "10010000",
1811 => "10010000",
1812 => "10010000",
1813 => "10010000",
1814 => "10010000",
1815 => "10010000",
1816 => "10010000",
1817 => "10010000",
1818 => "10010000",
1819 => "10010000",
1820 => "10010000",
1821 => "10010000",
1822 => "10010000",
1823 => "10010000",
1824 => "10010000",
1825 => "10010000",
1826 => "10010000",
1827 => "10010000",
1828 => "10010000",
1829 => "10010000",
1830 => "10010000",
1831 => "10010000",
1832 => "10010000",
1833 => "10010000",
1834 => "10010000",
1835 => "10010000",
1836 => "10010000",
1837 => "10010000",
1838 => "10010000",
1839 => "10010000",
1840 => "10010000",
1841 => "10010000",
1842 => "10010000",
1843 => "10010000",
1844 => "10010000",
1845 => "10010000",
1846 => "10010000",
1847 => "10010000",
1848 => "10010000",
1849 => "10010000",
1850 => "10010000",
1851 => "10010000",
1852 => "10010000",
1853 => "10010000",
1854 => "10010000",
1855 => "10010000",
1856 => "10010000",
1857 => "10010000",
1858 => "10010000",
1859 => "10010000",
1860 => "10010000",
1861 => "10010000",
1862 => "10010000",
1863 => "10010000",
1864 => "10010000",
1865 => "10010000",
1866 => "10010000",
1867 => "10010000",
1868 => "10010000",
1869 => "10010000",
1870 => "10010000",
1871 => "10010000",
1872 => "10010000",
1873 => "10010000",
1874 => "10010000",
1875 => "10010000",
1876 => "10010000",
1877 => "10010000",
1878 => "10010000",
1879 => "10010000",
1880 => "10010000",
1881 => "10010000",
1882 => "10010000",
1883 => "10010000",
1884 => "11111111",
1885 => "00000001",
1886 => "00000001",
1887 => "11111111",
1888 => "10010000",
1889 => "10010000",
1890 => "10010000",
1891 => "10010000",
1892 => "10010000",
1893 => "10010000",
1894 => "10010000",
1895 => "10010000",
1896 => "10010000",
1897 => "10010000",
1898 => "10010000",
1899 => "10010000",
1900 => "10010000",
1901 => "10010000",
1902 => "10010000",
1903 => "10010000",
1904 => "10010000",
1905 => "10010000",
1906 => "10010000",
1907 => "10010000",
1908 => "10010000",
1909 => "10010000",
1910 => "10010000",
1911 => "10010000",
1912 => "10010000",
1913 => "10010000",
1914 => "10010000",
1915 => "10010000",
1916 => "10010000",
1917 => "10010000",
1918 => "10010000",
1919 => "10010000",
1920 => "10010000",
1921 => "10010000",
1922 => "10010000",
1923 => "10010000",
1924 => "10010000",
1925 => "10010000",
1926 => "10010000",
1927 => "10010000",
1928 => "10010000",
1929 => "10010000",
1930 => "10010000",
1931 => "10010000",
1932 => "10010000",
1933 => "10010000",
1934 => "10010000",
1935 => "10010000",
1936 => "10010000",
1937 => "10010000",
1938 => "10010000",
1939 => "10010000",
1940 => "10010000",
1941 => "10010000",
1942 => "10010000",
1943 => "10010000",
1944 => "10010000",
1945 => "10010000",
1946 => "10010000",
1947 => "10010000",
1948 => "10010000",
1949 => "10010000",
1950 => "10010000",
1951 => "10010000",
1952 => "10010000",
1953 => "10010000",
1954 => "10010000",
1955 => "10010000",
1956 => "10010000",
1957 => "10010000",
1958 => "10010000",
1959 => "10010000",
1960 => "10010000",
1961 => "10010000",
1962 => "10010000",
1963 => "10010000",
1964 => "10010000",
1965 => "10010000",
1966 => "11111111",
1967 => "00000001",
1968 => "00000001",
1969 => "11111111",
1970 => "10010000",
1971 => "10010000",
1972 => "10010000",
1973 => "10010000",
1974 => "10010000",
1975 => "10010000",
1976 => "10010000",
1977 => "10010000",
1978 => "10010000",
1979 => "10010000",
1980 => "10010000",
1981 => "10010000",
1982 => "10010000",
1983 => "10010000",
1984 => "10010000",
1985 => "10010000",
1986 => "10010000",
1987 => "10010000",
1988 => "10010000",
1989 => "10010000",
1990 => "10010000",
1991 => "10010000",
1992 => "10010000",
1993 => "10010000",
1994 => "10010000",
1995 => "10010000",
1996 => "10010000",
1997 => "10010000",
1998 => "10010000",
1999 => "10010000",
2000 => "10010000",
2001 => "10010000",
2002 => "10010000",
2003 => "10010000",
2004 => "10010000",
2005 => "10010000",
2006 => "10010000",
2007 => "10010000",
2008 => "10010000",
2009 => "10010000",
2010 => "10010000",
2011 => "10010000",
2012 => "10010000",
2013 => "10010000",
2014 => "10010000",
2015 => "10010000",
2016 => "10010000",
2017 => "10010000",
2018 => "10010000",
2019 => "10010000",
2020 => "10010000",
2021 => "10010000",
2022 => "10010000",
2023 => "10010000",
2024 => "10010000",
2025 => "10010000",
2026 => "10010000",
2027 => "10010000",
2028 => "10010000",
2029 => "10010000",
2030 => "10010000",
2031 => "10010000",
2032 => "10010000",
2033 => "10010000",
2034 => "10010000",
2035 => "10010000",
2036 => "10010000",
2037 => "10010000",
2038 => "10010000",
2039 => "10010000",
2040 => "10010000",
2041 => "10010000",
2042 => "10010000",
2043 => "10010000",
2044 => "10010000",
2045 => "10010000",
2046 => "10010000",
2047 => "10010000",
2048 => "11111111",
2049 => "00000001",
2050 => "00000001",
2051 => "11111111",
2052 => "10010000",
2053 => "10010000",
2054 => "10010000",
2055 => "10010000",
2056 => "10010000",
2057 => "10010000",
2058 => "10010000",
2059 => "10010000",
2060 => "10010000",
2061 => "10010000",
2062 => "10010000",
2063 => "10010000",
2064 => "10010000",
2065 => "10010000",
2066 => "10010000",
2067 => "10010000",
2068 => "10010000",
2069 => "10010000",
2070 => "10010000",
2071 => "10010000",
2072 => "10010000",
2073 => "10010000",
2074 => "10010000",
2075 => "10010000",
2076 => "10010000",
2077 => "10010000",
2078 => "10010000",
2079 => "10010000",
2080 => "10010000",
2081 => "10010000",
2082 => "10010000",
2083 => "10010000",
2084 => "10010000",
2085 => "10010000",
2086 => "10010000",
2087 => "10010000",
2088 => "10010000",
2089 => "10010000",
2090 => "10010000",
2091 => "10010000",
2092 => "10010000",
2093 => "10010000",
2094 => "10010000",
2095 => "10010000",
2096 => "10010000",
2097 => "10010000",
2098 => "10010000",
2099 => "10010000",
2100 => "10010000",
2101 => "10010000",
2102 => "10010000",
2103 => "10010000",
2104 => "10010000",
2105 => "10010000",
2106 => "10010000",
2107 => "10010000",
2108 => "10010000",
2109 => "10010000",
2110 => "10010000",
2111 => "10010000",
2112 => "10010000",
2113 => "10010000",
2114 => "10010000",
2115 => "10010000",
2116 => "10010000",
2117 => "10010000",
2118 => "10010000",
2119 => "10010000",
2120 => "10010000",
2121 => "10010000",
2122 => "10010000",
2123 => "10010000",
2124 => "10010000",
2125 => "10010000",
2126 => "10010000",
2127 => "10010000",
2128 => "10010000",
2129 => "10010000",
2130 => "11111111",
2131 => "00000001",
2132 => "00000001",
2133 => "11111111",
2134 => "10010000",
2135 => "10010000",
2136 => "10010000",
2137 => "10010000",
2138 => "10010000",
2139 => "10010000",
2140 => "10010000",
2141 => "10010000",
2142 => "10010000",
2143 => "10010000",
2144 => "10010000",
2145 => "10010000",
2146 => "10010000",
2147 => "10010000",
2148 => "10010000",
2149 => "10010000",
2150 => "10010000",
2151 => "10010000",
2152 => "10010000",
2153 => "10010000",
2154 => "10010000",
2155 => "10010000",
2156 => "10010000",
2157 => "10010000",
2158 => "10010000",
2159 => "10010000",
2160 => "10010000",
2161 => "10010000",
2162 => "10010000",
2163 => "10010000",
2164 => "10010000",
2165 => "10010000",
2166 => "10010000",
2167 => "10010000",
2168 => "10010000",
2169 => "10010000",
2170 => "10010000",
2171 => "10010000",
2172 => "10010000",
2173 => "10010000",
2174 => "10010000",
2175 => "10010000",
2176 => "10010000",
2177 => "10010000",
2178 => "10010000",
2179 => "10010000",
2180 => "10010000",
2181 => "10010000",
2182 => "10010000",
2183 => "10010000",
2184 => "10010000",
2185 => "10010000",
2186 => "10010000",
2187 => "10010000",
2188 => "10010000",
2189 => "10010000",
2190 => "10010000",
2191 => "10010000",
2192 => "10010000",
2193 => "10010000",
2194 => "10010000",
2195 => "10010000",
2196 => "10010000",
2197 => "10010000",
2198 => "10010000",
2199 => "10010000",
2200 => "10010000",
2201 => "10010000",
2202 => "10010000",
2203 => "10010000",
2204 => "10010000",
2205 => "10010000",
2206 => "10010000",
2207 => "10010000",
2208 => "10010000",
2209 => "10010000",
2210 => "10010000",
2211 => "10010000",
2212 => "11111111",
2213 => "00000001",
2214 => "00000001",
2215 => "11111111",
2216 => "10010000",
2217 => "10010000",
2218 => "10010000",
2219 => "10010000",
2220 => "10010000",
2221 => "10010000",
2222 => "10010000",
2223 => "10010000",
2224 => "10010000",
2225 => "10010000",
2226 => "10010000",
2227 => "10010000",
2228 => "10010000",
2229 => "10010000",
2230 => "10010000",
2231 => "10010000",
2232 => "10010000",
2233 => "10010000",
2234 => "10010000",
2235 => "10010000",
2236 => "10010000",
2237 => "10010000",
2238 => "10010000",
2239 => "10010000",
2240 => "10010000",
2241 => "10010000",
2242 => "10010000",
2243 => "10010000",
2244 => "10010000",
2245 => "10010000",
2246 => "10010000",
2247 => "10010000",
2248 => "10010000",
2249 => "10010000",
2250 => "10010000",
2251 => "10010000",
2252 => "10010000",
2253 => "10010000",
2254 => "10010000",
2255 => "10010000",
2256 => "10010000",
2257 => "10010000",
2258 => "10010000",
2259 => "10010000",
2260 => "10010000",
2261 => "10010000",
2262 => "10010000",
2263 => "10010000",
2264 => "10010000",
2265 => "10010000",
2266 => "10010000",
2267 => "10010000",
2268 => "10010000",
2269 => "10010000",
2270 => "10010000",
2271 => "10010000",
2272 => "10010000",
2273 => "10010000",
2274 => "10010000",
2275 => "10010000",
2276 => "10010000",
2277 => "10010000",
2278 => "10010000",
2279 => "10010000",
2280 => "10010000",
2281 => "10010000",
2282 => "10010000",
2283 => "10010000",
2284 => "10010000",
2285 => "10010000",
2286 => "10010000",
2287 => "10010000",
2288 => "10010000",
2289 => "10010000",
2290 => "10010000",
2291 => "10010000",
2292 => "10010000",
2293 => "10010000",
2294 => "11111111",
2295 => "00000001",
2296 => "00000001",
2297 => "10110110",
2298 => "10110101",
2299 => "10010000",
2300 => "10010000",
2301 => "10010000",
2302 => "10010000",
2303 => "10010000",
2304 => "10010000",
2305 => "10010000",
2306 => "10010000",
2307 => "10010000",
2308 => "10010000",
2309 => "10010000",
2310 => "10010000",
2311 => "10010000",
2312 => "10010000",
2313 => "10010000",
2314 => "10010000",
2315 => "10010000",
2316 => "10010000",
2317 => "10010000",
2318 => "10010000",
2319 => "10010000",
2320 => "10010000",
2321 => "10010000",
2322 => "10010000",
2323 => "10010000",
2324 => "10010000",
2325 => "10010000",
2326 => "10010000",
2327 => "10010000",
2328 => "10010000",
2329 => "10010000",
2330 => "10010000",
2331 => "10010000",
2332 => "10010000",
2333 => "10010000",
2334 => "10010000",
2335 => "10010000",
2336 => "10010000",
2337 => "10010000",
2338 => "10010000",
2339 => "10010000",
2340 => "10010000",
2341 => "10010000",
2342 => "10010000",
2343 => "10010000",
2344 => "10010000",
2345 => "10010000",
2346 => "10010000",
2347 => "10010000",
2348 => "10010000",
2349 => "10010000",
2350 => "10010000",
2351 => "10010000",
2352 => "10010000",
2353 => "10010000",
2354 => "10010000",
2355 => "10010000",
2356 => "10010000",
2357 => "10010000",
2358 => "10010000",
2359 => "10010000",
2360 => "10010000",
2361 => "10010000",
2362 => "10010000",
2363 => "10010000",
2364 => "10010000",
2365 => "10010000",
2366 => "10010000",
2367 => "10010000",
2368 => "10010000",
2369 => "10010000",
2370 => "10010000",
2371 => "10010000",
2372 => "10010000",
2373 => "10010000",
2374 => "10010000",
2375 => "10110101",
2376 => "10110110",
2377 => "00000001",
2378 => "00000001",
2379 => "00100101",
2380 => "11111111",
2381 => "10110101",
2382 => "10010000",
2383 => "10010000",
2384 => "10010000",
2385 => "10010000",
2386 => "10010000",
2387 => "10010000",
2388 => "10010000",
2389 => "10010000",
2390 => "10010000",
2391 => "10010000",
2392 => "10010000",
2393 => "10010000",
2394 => "10010000",
2395 => "10010000",
2396 => "10010000",
2397 => "10010000",
2398 => "10010000",
2399 => "10010000",
2400 => "10010000",
2401 => "10010000",
2402 => "10010000",
2403 => "10010000",
2404 => "10010000",
2405 => "10010000",
2406 => "10010000",
2407 => "10010000",
2408 => "10010000",
2409 => "10010000",
2410 => "10010000",
2411 => "10010000",
2412 => "10010000",
2413 => "10010000",
2414 => "10010000",
2415 => "10010000",
2416 => "10010000",
2417 => "10010000",
2418 => "10010000",
2419 => "10010000",
2420 => "10010000",
2421 => "10010000",
2422 => "10010000",
2423 => "10010000",
2424 => "10010000",
2425 => "10010000",
2426 => "10010000",
2427 => "10010000",
2428 => "10010000",
2429 => "10010000",
2430 => "10010000",
2431 => "10010000",
2432 => "10010000",
2433 => "10010000",
2434 => "10010000",
2435 => "10010000",
2436 => "10010000",
2437 => "10010000",
2438 => "10010000",
2439 => "10010000",
2440 => "10010000",
2441 => "10010000",
2442 => "10010000",
2443 => "10010000",
2444 => "10010000",
2445 => "10010000",
2446 => "10010000",
2447 => "10010000",
2448 => "10010000",
2449 => "10010000",
2450 => "10010000",
2451 => "10010000",
2452 => "10010000",
2453 => "10010000",
2454 => "10010000",
2455 => "10010000",
2456 => "10110101",
2457 => "11111111",
2458 => "00100101",
2459 => "00000001",
2460 => "00000001",
2461 => "00000001",
2462 => "00100101",
2463 => "10110110",
2464 => "11111111",
2465 => "11111111",
2466 => "11111111",
2467 => "11111111",
2468 => "11111111",
2469 => "11111111",
2470 => "11111111",
2471 => "11111111",
2472 => "11111111",
2473 => "11111111",
2474 => "11111111",
2475 => "11111111",
2476 => "11111111",
2477 => "11111111",
2478 => "11111111",
2479 => "11111111",
2480 => "11111111",
2481 => "11111111",
2482 => "11111111",
2483 => "11111111",
2484 => "11111111",
2485 => "11111111",
2486 => "11111111",
2487 => "11111111",
2488 => "11111111",
2489 => "11111111",
2490 => "11111111",
2491 => "11111111",
2492 => "11111111",
2493 => "11111111",
2494 => "11111111",
2495 => "11111111",
2496 => "11111111",
2497 => "11111111",
2498 => "11111111",
2499 => "11111111",
2500 => "11111111",
2501 => "11111111",
2502 => "11111111",
2503 => "11111111",
2504 => "11111111",
2505 => "11111111",
2506 => "11111111",
2507 => "11111111",
2508 => "11111111",
2509 => "11111111",
2510 => "11111111",
2511 => "11111111",
2512 => "11111111",
2513 => "11111111",
2514 => "11111111",
2515 => "11111111",
2516 => "11111111",
2517 => "11111111",
2518 => "11111111",
2519 => "11111111",
2520 => "11111111",
2521 => "11111111",
2522 => "11111111",
2523 => "11111111",
2524 => "11111111",
2525 => "11111111",
2526 => "11111111",
2527 => "11111111",
2528 => "11111111",
2529 => "11111111",
2530 => "11111111",
2531 => "11111111",
2532 => "11111111",
2533 => "11111111",
2534 => "11111111",
2535 => "11111111",
2536 => "11111111",
2537 => "11111111",
2538 => "10110110",
2539 => "00100101",
2540 => "00000001",
2541 => "00000001",
2542 => "00000001",
2543 => "00000001",
2544 => "00000001",
2545 => "00000001",
2546 => "00000001",
2547 => "00000001",
2548 => "00000001",
2549 => "00000001",
2550 => "00000001",
2551 => "00000001",
2552 => "00000001",
2553 => "00000001",
2554 => "00000001",
2555 => "00000001",
2556 => "00000001",
2557 => "00000001",
2558 => "00000001",
2559 => "00000001",
2560 => "00000001",
2561 => "00000001",
2562 => "00000001",
2563 => "00000001",
2564 => "00000001",
2565 => "00000001",
2566 => "00000001",
2567 => "00000001",
2568 => "00000001",
2569 => "00000001",
2570 => "00000001",
2571 => "00000001",
2572 => "00000001",
2573 => "00000001",
2574 => "00000001",
2575 => "00000001",
2576 => "00000001",
2577 => "00000001",
2578 => "00000001",
2579 => "00000001",
2580 => "00000001",
2581 => "00000001",
2582 => "00000001",
2583 => "00000001",
2584 => "00000001",
2585 => "00000001",
2586 => "00000001",
2587 => "00000001",
2588 => "00000001",
2589 => "00000001",
2590 => "00000001",
2591 => "00000001",
2592 => "00000001",
2593 => "00000001",
2594 => "00000001",
2595 => "00000001",
2596 => "00000001",
2597 => "00000001",
2598 => "00000001",
2599 => "00000001",
2600 => "00000001",
2601 => "00000001",
2602 => "00000001",
2603 => "00000001",
2604 => "00000001",
2605 => "00000001",
2606 => "00000001",
2607 => "00000001",
2608 => "00000001",
2609 => "00000001",
2610 => "00000001",
2611 => "00000001",
2612 => "00000001",
2613 => "00000001",
2614 => "00000001",
2615 => "00000001",
2616 => "00000001",
2617 => "00000001",
2618 => "00000001",
2619 => "00000001",
2620 => "00000001",
2621 => "00000001",
2622 => "00000001",
2623 => "00000001");
begin

    process(clk)
    begin
    
        if rising_edge(clk) then
                dout <= yellow(to_integer(unsigned(addr)));
        end if;
    end process;

end Behavioral;

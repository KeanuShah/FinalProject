
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity Button_Live is
    port(clk, rst: in std_logic;
         addr: in std_logic_vector(11 downto 0);
         dout: out std_logic_vector(7 downto 0));
end Button_Live;

architecture Behavioral of Button_Live is

 type mem is array (0 to 2749) of std_logic_vector(7 downto 0);
 signal live: mem:= (
    0 => "00000001",
        1 => "00000001",
        2 => "00000001",
        3 => "00000001",
        4 => "00000001",
        5 => "00000001",
        6 => "00000001",
        7 => "00000001",
        8 => "00000001",
        9 => "00000001",
        10 => "00000001",
        11 => "00000001",
        12 => "00000001",
        13 => "00000001",
        14 => "00000001",
        15 => "00000001",
        16 => "00000001",
        17 => "00000001",
        18 => "00000001",
        19 => "00000001",
        20 => "00000001",
        21 => "00000001",
        22 => "00000001",
        23 => "00000001",
        24 => "00000001",
        25 => "00000001",
        26 => "00000001",
        27 => "00000001",
        28 => "00000001",
        29 => "00000001",
        30 => "00000001",
        31 => "00000001",
        32 => "00000001",
        33 => "00000001",
        34 => "00000001",
        35 => "00000001",
        36 => "00000001",
        37 => "00000001",
        38 => "00000001",
        39 => "00000001",
        40 => "00000001",
        41 => "00000001",
        42 => "00000001",
        43 => "00000001",
        44 => "00000001",
        45 => "00000001",
        46 => "00000001",
        47 => "00000001",
        48 => "00000001",
        49 => "00000001",
        50 => "00000001",
        51 => "00000001",
        52 => "00000001",
        53 => "00000001",
        54 => "00000001",
        55 => "00000001",
        56 => "00000001",
        57 => "00000001",
        58 => "00000001",
        59 => "00000001",
        60 => "00000001",
        61 => "00000001",
        62 => "00000001",
        63 => "00000001",
        64 => "00000001",
        65 => "00000001",
        66 => "00000001",
        67 => "00000001",
        68 => "00000001",
        69 => "00000001",
        70 => "00000001",
        71 => "00000001",
        72 => "00000001",
        73 => "00000001",
        74 => "00000001",
        75 => "00000001",
        76 => "00000001",
        77 => "00000001",
        78 => "00000001",
        79 => "00000001",
        80 => "00000001",
        81 => "00000001",
        82 => "00000001",
        83 => "00000001",
        84 => "00000001",
        85 => "00000001",
        86 => "00000001",
        87 => "00000001",
        88 => "00000001",
        89 => "00000001",
        90 => "00000001",
        91 => "00000001",
        92 => "00000001",
        93 => "00000001",
        94 => "00000001",
        95 => "00000001",
        96 => "00000001",
        97 => "00000001",
        98 => "00000001",
        99 => "00000001",
        100 => "00000001",
        101 => "00000001",
        102 => "00000001",
        103 => "00000001",
        104 => "00000001",
        105 => "00000001",
        106 => "00000001",
        107 => "00000001",
        108 => "00000001",
        109 => "00000001",
        110 => "00000001",
        111 => "00000001",
        112 => "00100101",
        113 => "10110110",
        114 => "11111111",
        115 => "11111111",
        116 => "11111111",
        117 => "11111111",
        118 => "11111111",
        119 => "11111111",
        120 => "11111111",
        121 => "11111111",
        122 => "11111111",
        123 => "11111111",
        124 => "11111111",
        125 => "11111111",
        126 => "11111111",
        127 => "11111111",
        128 => "11111111",
        129 => "11111111",
        130 => "11111111",
        131 => "11111111",
        132 => "11111111",
        133 => "11111111",
        134 => "11111111",
        135 => "11111111",
        136 => "11111111",
        137 => "11111111",
        138 => "11111111",
        139 => "11111111",
        140 => "11111111",
        141 => "11111111",
        142 => "11111111",
        143 => "11111111",
        144 => "11111111",
        145 => "11111111",
        146 => "11111111",
        147 => "11111111",
        148 => "11111111",
        149 => "11111111",
        150 => "11111111",
        151 => "11111111",
        152 => "11111111",
        153 => "11111111",
        154 => "11111111",
        155 => "11111111",
        156 => "11111111",
        157 => "11111111",
        158 => "11111111",
        159 => "11111111",
        160 => "11111111",
        161 => "11111111",
        162 => "11111111",
        163 => "11111111",
        164 => "11111111",
        165 => "11111111",
        166 => "11111111",
        167 => "11111111",
        168 => "11111111",
        169 => "11111111",
        170 => "11111111",
        171 => "11111111",
        172 => "11111111",
        173 => "11111111",
        174 => "11111111",
        175 => "11111111",
        176 => "11111111",
        177 => "11111111",
        178 => "11111111",
        179 => "11111111",
        180 => "11111111",
        181 => "11111111",
        182 => "11111111",
        183 => "11111111",
        184 => "11111111",
        185 => "11111111",
        186 => "11111111",
        187 => "11111111",
        188 => "11111111",
        189 => "11111111",
        190 => "11111111",
        191 => "11111111",
        192 => "11111111",
        193 => "11111111",
        194 => "11111111",
        195 => "11111111",
        196 => "11111111",
        197 => "11111111",
        198 => "11111111",
        199 => "11111111",
        200 => "11111111",
        201 => "11111111",
        202 => "11111111",
        203 => "11111111",
        204 => "11111111",
        205 => "11111111",
        206 => "11111111",
        207 => "11111111",
        208 => "11111111",
        209 => "11111111",
        210 => "11111111",
        211 => "11111111",
        212 => "11111111",
        213 => "11111111",
        214 => "11111111",
        215 => "11111111",
        216 => "10110110",
        217 => "00100101",
        218 => "00000001",
        219 => "00000001",
        220 => "00000001",
        221 => "00100101",
        222 => "11111111",
        223 => "11111111",
        224 => "11111111",
        225 => "11111111",
        226 => "11111111",
        227 => "11111111",
        228 => "11111111",
        229 => "11111111",
        230 => "11111111",
        231 => "11111111",
        232 => "11111111",
        233 => "11111111",
        234 => "11111111",
        235 => "11111111",
        236 => "11111111",
        237 => "11111111",
        238 => "11111111",
        239 => "11111111",
        240 => "11111111",
        241 => "11111111",
        242 => "11111111",
        243 => "11111111",
        244 => "11111111",
        245 => "11111111",
        246 => "11111111",
        247 => "11111111",
        248 => "11111111",
        249 => "11111111",
        250 => "11111111",
        251 => "11111111",
        252 => "11111111",
        253 => "11111111",
        254 => "11111111",
        255 => "11111111",
        256 => "11111111",
        257 => "11111111",
        258 => "11111111",
        259 => "11111111",
        260 => "11111111",
        261 => "11111111",
        262 => "11111111",
        263 => "11111111",
        264 => "11111111",
        265 => "11111111",
        266 => "11111111",
        267 => "11111111",
        268 => "11111111",
        269 => "11111111",
        270 => "11111111",
        271 => "11111111",
        272 => "11111111",
        273 => "11111111",
        274 => "11111111",
        275 => "11111111",
        276 => "11111111",
        277 => "11111111",
        278 => "11111111",
        279 => "11111111",
        280 => "11111111",
        281 => "11111111",
        282 => "11111111",
        283 => "11111111",
        284 => "11111111",
        285 => "11111111",
        286 => "11111111",
        287 => "11111111",
        288 => "11111111",
        289 => "11111111",
        290 => "11111111",
        291 => "11111111",
        292 => "11111111",
        293 => "11111111",
        294 => "11111111",
        295 => "11111111",
        296 => "11111111",
        297 => "11111111",
        298 => "11111111",
        299 => "11111111",
        300 => "11111111",
        301 => "11111111",
        302 => "11111111",
        303 => "11111111",
        304 => "11111111",
        305 => "11111111",
        306 => "11111111",
        307 => "11111111",
        308 => "11111111",
        309 => "11111111",
        310 => "11111111",
        311 => "11111111",
        312 => "11111111",
        313 => "11111111",
        314 => "11111111",
        315 => "11111111",
        316 => "11111111",
        317 => "11111111",
        318 => "11111111",
        319 => "11111111",
        320 => "11111111",
        321 => "11111111",
        322 => "11111111",
        323 => "11111111",
        324 => "11111111",
        325 => "11111111",
        326 => "11111111",
        327 => "11111111",
        328 => "00100101",
        329 => "00000001",
        330 => "00000001",
        331 => "10110110",
        332 => "11111111",
        333 => "01010001",
        334 => "00010100",
        335 => "00010100",
        336 => "00010100",
        337 => "00010100",
        338 => "00010100",
        339 => "00010100",
        340 => "00010100",
        341 => "00010100",
        342 => "00010100",
        343 => "00010100",
        344 => "00010100",
        345 => "00010100",
        346 => "00010100",
        347 => "00010100",
        348 => "00010100",
        349 => "00010100",
        350 => "00010100",
        351 => "00010100",
        352 => "00010100",
        353 => "00010100",
        354 => "00010100",
        355 => "00010100",
        356 => "00010100",
        357 => "00010100",
        358 => "00010100",
        359 => "00010100",
        360 => "00010100",
        361 => "00010100",
        362 => "00010100",
        363 => "00010100",
        364 => "00010100",
        365 => "00010100",
        366 => "00010100",
        367 => "00010100",
        368 => "00010100",
        369 => "00010100",
        370 => "00010100",
        371 => "00010100",
        372 => "00010100",
        373 => "00010100",
        374 => "00010100",
        375 => "00010100",
        376 => "00010100",
        377 => "00010100",
        378 => "00010100",
        379 => "00010100",
        380 => "00010100",
        381 => "00010100",
        382 => "00010100",
        383 => "00010100",
        384 => "00010100",
        385 => "00000001",
        386 => "00000001",
        387 => "00000001",
        388 => "00000001",
        389 => "00000001",
        390 => "00000001",
        391 => "00000001",
        392 => "00000001",
        393 => "00000001",
        394 => "00000001",
        395 => "00000001",
        396 => "00000001",
        397 => "00000001",
        398 => "00000001",
        399 => "00000001",
        400 => "00000001",
        401 => "00000001",
        402 => "00000001",
        403 => "00000001",
        404 => "00000001",
        405 => "00000001",
        406 => "00000001",
        407 => "00000001",
        408 => "00000001",
        409 => "00000001",
        410 => "00000001",
        411 => "00000001",
        412 => "00000001",
        413 => "00000001",
        414 => "00000001",
        415 => "00000001",
        416 => "00000001",
        417 => "00000001",
        418 => "00000001",
        419 => "00000001",
        420 => "00000001",
        421 => "00000001",
        422 => "00000001",
        423 => "00000001",
        424 => "00000001",
        425 => "00000001",
        426 => "00000001",
        427 => "00000001",
        428 => "00000001",
        429 => "00000001",
        430 => "00000001",
        431 => "00000001",
        432 => "00000001",
        433 => "00000001",
        434 => "00000001",
        435 => "00000001",
        436 => "01001010",
        437 => "11111111",
        438 => "10110110",
        439 => "00000001",
        440 => "00000001",
        441 => "11111111",
        442 => "11111111",
        443 => "00010100",
        444 => "00010100",
        445 => "00010100",
        446 => "00010100",
        447 => "00010100",
        448 => "00010100",
        449 => "00010100",
        450 => "00010100",
        451 => "00010100",
        452 => "00010100",
        453 => "00010100",
        454 => "00010100",
        455 => "00010100",
        456 => "00010100",
        457 => "00010100",
        458 => "00010100",
        459 => "00010100",
        460 => "00010100",
        461 => "00010100",
        462 => "00010100",
        463 => "00010100",
        464 => "00010100",
        465 => "00010100",
        466 => "00010100",
        467 => "00010100",
        468 => "00010100",
        469 => "00010100",
        470 => "00010100",
        471 => "00010100",
        472 => "00010100",
        473 => "00010100",
        474 => "00010100",
        475 => "00010100",
        476 => "00010100",
        477 => "00010100",
        478 => "00010100",
        479 => "00010100",
        480 => "00010100",
        481 => "00010100",
        482 => "00010100",
        483 => "00010100",
        484 => "00010100",
        485 => "00010100",
        486 => "00010100",
        487 => "00010100",
        488 => "00010100",
        489 => "00010100",
        490 => "00010100",
        491 => "00010100",
        492 => "00010100",
        493 => "00010100",
        494 => "00010100",
        495 => "00000001",
        496 => "00000001",
        497 => "00000001",
        498 => "00000001",
        499 => "00000001",
        500 => "00000001",
        501 => "00000001",
        502 => "00000001",
        503 => "00000001",
        504 => "00000001",
        505 => "00000001",
        506 => "00000001",
        507 => "00000001",
        508 => "00000001",
        509 => "00000001",
        510 => "00000001",
        511 => "00000001",
        512 => "00000001",
        513 => "00000001",
        514 => "00000001",
        515 => "00000001",
        516 => "00000001",
        517 => "00000001",
        518 => "00000001",
        519 => "00000001",
        520 => "00000001",
        521 => "00000001",
        522 => "00000001",
        523 => "00000001",
        524 => "00000001",
        525 => "00000001",
        526 => "00000001",
        527 => "00000001",
        528 => "00000001",
        529 => "00000001",
        530 => "00000001",
        531 => "00000001",
        532 => "00000001",
        533 => "00000001",
        534 => "00000001",
        535 => "00000001",
        536 => "00000001",
        537 => "00000001",
        538 => "00000001",
        539 => "00000001",
        540 => "00000001",
        541 => "00000001",
        542 => "00000001",
        543 => "00000001",
        544 => "00000001",
        545 => "00000001",
        546 => "00000001",
        547 => "11111111",
        548 => "11111111",
        549 => "00000001",
        550 => "00000001",
        551 => "11111111",
        552 => "11111111",
        553 => "00010100",
        554 => "00010100",
        555 => "00010100",
        556 => "00010100",
        557 => "00010100",
        558 => "00010100",
        559 => "00010100",
        560 => "00010100",
        561 => "00010100",
        562 => "00010100",
        563 => "00010100",
        564 => "00010100",
        565 => "00010100",
        566 => "00010100",
        567 => "00010100",
        568 => "00010100",
        569 => "00010100",
        570 => "00010100",
        571 => "00010100",
        572 => "00010100",
        573 => "00010100",
        574 => "00010100",
        575 => "00010100",
        576 => "00010100",
        577 => "00010100",
        578 => "00010100",
        579 => "00010100",
        580 => "00010100",
        581 => "00010100",
        582 => "00010100",
        583 => "00010100",
        584 => "00010100",
        585 => "00010100",
        586 => "00010100",
        587 => "00010100",
        588 => "00010100",
        589 => "00010100",
        590 => "00010100",
        591 => "00010100",
        592 => "00010100",
        593 => "00010100",
        594 => "00010100",
        595 => "00010100",
        596 => "00010100",
        597 => "00010100",
        598 => "00010100",
        599 => "00010100",
        600 => "00010100",
        601 => "00010100",
        602 => "00010100",
        603 => "00010100",
        604 => "00010100",
        605 => "00000001",
        606 => "00000001",
        607 => "00000001",
        608 => "00000001",
        609 => "00000001",
        610 => "00000001",
        611 => "00000001",
        612 => "00000001",
        613 => "00000001",
        614 => "00000001",
        615 => "00000001",
        616 => "00000001",
        617 => "00000001",
        618 => "00000001",
        619 => "00000001",
        620 => "00000001",
        621 => "00000001",
        622 => "00000001",
        623 => "00000001",
        624 => "00000001",
        625 => "00000001",
        626 => "00000001",
        627 => "00000001",
        628 => "00000001",
        629 => "00000001",
        630 => "00000001",
        631 => "00000001",
        632 => "00000001",
        633 => "00000001",
        634 => "00000001",
        635 => "00000001",
        636 => "00000001",
        637 => "00000001",
        638 => "00000001",
        639 => "00000001",
        640 => "00000001",
        641 => "00000001",
        642 => "00000001",
        643 => "00000001",
        644 => "00000001",
        645 => "00000001",
        646 => "00000001",
        647 => "00000001",
        648 => "00000001",
        649 => "00000001",
        650 => "00000001",
        651 => "00000001",
        652 => "00000001",
        653 => "00000001",
        654 => "00000001",
        655 => "00000001",
        656 => "00000001",
        657 => "11111111",
        658 => "11111111",
        659 => "00000001",
        660 => "00000001",
        661 => "11111111",
        662 => "11111111",
        663 => "00010100",
        664 => "00010100",
        665 => "00010100",
        666 => "00010100",
        667 => "00010100",
        668 => "00010100",
        669 => "00010100",
        670 => "00010100",
        671 => "00010100",
        672 => "00010100",
        673 => "00010100",
        674 => "00010100",
        675 => "00010100",
        676 => "00010100",
        677 => "00010100",
        678 => "00010100",
        679 => "00010100",
        680 => "00010100",
        681 => "00010100",
        682 => "00010100",
        683 => "00010100",
        684 => "00010100",
        685 => "00010100",
        686 => "00010100",
        687 => "00010100",
        688 => "00010100",
        689 => "00010100",
        690 => "00010100",
        691 => "00010100",
        692 => "00010100",
        693 => "00010100",
        694 => "00010100",
        695 => "00010100",
        696 => "00010100",
        697 => "00010100",
        698 => "00010100",
        699 => "00010100",
        700 => "00010100",
        701 => "00010100",
        702 => "00010100",
        703 => "00010100",
        704 => "00010100",
        705 => "00010100",
        706 => "00010100",
        707 => "00010100",
        708 => "00010100",
        709 => "00010100",
        710 => "00010100",
        711 => "00010100",
        712 => "00010100",
        713 => "00010100",
        714 => "00010100",
        715 => "00000001",
        716 => "00000001",
        717 => "00000001",
        718 => "00000001",
        719 => "00000001",
        720 => "00000001",
        721 => "00000001",
        722 => "00000001",
        723 => "00000001",
        724 => "00000001",
        725 => "00000001",
        726 => "00000001",
        727 => "00000001",
        728 => "00000001",
        729 => "00000001",
        730 => "00000001",
        731 => "00000001",
        732 => "00000001",
        733 => "00000001",
        734 => "00000001",
        735 => "00000001",
        736 => "00000001",
        737 => "00000001",
        738 => "00000001",
        739 => "00000001",
        740 => "00000001",
        741 => "00000001",
        742 => "00000001",
        743 => "00000001",
        744 => "00000001",
        745 => "00000001",
        746 => "00000001",
        747 => "00000001",
        748 => "00000001",
        749 => "00000001",
        750 => "00000001",
        751 => "00000001",
        752 => "00000001",
        753 => "00000001",
        754 => "00000001",
        755 => "00000001",
        756 => "00000001",
        757 => "00000001",
        758 => "00000001",
        759 => "00000001",
        760 => "00000001",
        761 => "00000001",
        762 => "00000001",
        763 => "00000001",
        764 => "00000001",
        765 => "00000001",
        766 => "00000001",
        767 => "11111111",
        768 => "11111111",
        769 => "00000001",
        770 => "00000001",
        771 => "11111111",
        772 => "11111111",
        773 => "00010100",
        774 => "00010100",
        775 => "00010100",
        776 => "00010100",
        777 => "00010100",
        778 => "00010100",
        779 => "00010100",
        780 => "00010100",
        781 => "00010100",
        782 => "00010100",
        783 => "00010100",
        784 => "00010100",
        785 => "00010100",
        786 => "00010100",
        787 => "00010100",
        788 => "00010100",
        789 => "00010100",
        790 => "00010100",
        791 => "00010100",
        792 => "00010100",
        793 => "00010100",
        794 => "00010100",
        795 => "00010100",
        796 => "00010100",
        797 => "00010100",
        798 => "00010100",
        799 => "00010100",
        800 => "00010100",
        801 => "00010100",
        802 => "00010100",
        803 => "00010100",
        804 => "00010100",
        805 => "00010100",
        806 => "00010100",
        807 => "00010100",
        808 => "00010100",
        809 => "00010100",
        810 => "00010100",
        811 => "00010100",
        812 => "00010100",
        813 => "00010100",
        814 => "00010100",
        815 => "00010100",
        816 => "00010100",
        817 => "00010100",
        818 => "00010100",
        819 => "00010100",
        820 => "00010100",
        821 => "00010100",
        822 => "00010100",
        823 => "00010100",
        824 => "00010100",
        825 => "00000001",
        826 => "00000001",
        827 => "00000001",
        828 => "00000001",
        829 => "00000001",
        830 => "00000001",
        831 => "00000001",
        832 => "00000001",
        833 => "00000001",
        834 => "00000001",
        835 => "00000001",
        836 => "00000001",
        837 => "00000001",
        838 => "00000001",
        839 => "00000001",
        840 => "00000001",
        841 => "00000001",
        842 => "00000001",
        843 => "00000001",
        844 => "00000001",
        845 => "00000001",
        846 => "00000001",
        847 => "00000001",
        848 => "00000001",
        849 => "00000001",
        850 => "00000001",
        851 => "00000001",
        852 => "00000001",
        853 => "00000001",
        854 => "00000001",
        855 => "00000001",
        856 => "00000001",
        857 => "00000001",
        858 => "00000001",
        859 => "00000001",
        860 => "00000001",
        861 => "00000001",
        862 => "00000001",
        863 => "00000001",
        864 => "00000001",
        865 => "00000001",
        866 => "00000001",
        867 => "00000001",
        868 => "00000001",
        869 => "00000001",
        870 => "00000001",
        871 => "00000001",
        872 => "00000001",
        873 => "00000001",
        874 => "00000001",
        875 => "00000001",
        876 => "00000001",
        877 => "11111111",
        878 => "11111111",
        879 => "00000001",
        880 => "00000001",
        881 => "11111111",
        882 => "11111111",
        883 => "00010100",
        884 => "00010100",
        885 => "00010100",
        886 => "00010100",
        887 => "00010100",
        888 => "00010100",
        889 => "00010100",
        890 => "00010100",
        891 => "00010100",
        892 => "00010100",
        893 => "00010100",
        894 => "00010100",
        895 => "00010100",
        896 => "00010100",
        897 => "00010100",
        898 => "00010100",
        899 => "00010100",
        900 => "00010100",
        901 => "00010100",
        902 => "00010100",
        903 => "00010100",
        904 => "00010100",
        905 => "00010100",
        906 => "00010100",
        907 => "00010100",
        908 => "00010100",
        909 => "00010100",
        910 => "00010100",
        911 => "00010100",
        912 => "00010100",
        913 => "00010100",
        914 => "00010100",
        915 => "00010100",
        916 => "00010100",
        917 => "00010100",
        918 => "00010100",
        919 => "00010100",
        920 => "00010100",
        921 => "00010100",
        922 => "00010100",
        923 => "00010100",
        924 => "00010100",
        925 => "00010100",
        926 => "00010100",
        927 => "00010100",
        928 => "00010100",
        929 => "00010100",
        930 => "00010100",
        931 => "00010100",
        932 => "00010100",
        933 => "00010100",
        934 => "00010100",
        935 => "00000001",
        936 => "00000001",
        937 => "00000001",
        938 => "00000001",
        939 => "00000001",
        940 => "00000001",
        941 => "00000001",
        942 => "00000001",
        943 => "00000001",
        944 => "00000001",
        945 => "00000001",
        946 => "00000001",
        947 => "00000001",
        948 => "00000001",
        949 => "00000001",
        950 => "00000001",
        951 => "00000001",
        952 => "00000001",
        953 => "00000001",
        954 => "00000001",
        955 => "00000001",
        956 => "00000001",
        957 => "00000001",
        958 => "00000001",
        959 => "00000001",
        960 => "00000001",
        961 => "00000001",
        962 => "00000001",
        963 => "00000001",
        964 => "00000001",
        965 => "00000001",
        966 => "00000001",
        967 => "00000001",
        968 => "00000001",
        969 => "00000001",
        970 => "00000001",
        971 => "00000001",
        972 => "00000001",
        973 => "00000001",
        974 => "00000001",
        975 => "00000001",
        976 => "00000001",
        977 => "00000001",
        978 => "00000001",
        979 => "00000001",
        980 => "00000001",
        981 => "00000001",
        982 => "00000001",
        983 => "00000001",
        984 => "00000001",
        985 => "00000001",
        986 => "00000001",
        987 => "11111111",
        988 => "11111111",
        989 => "00000001",
        990 => "00000001",
        991 => "11111111",
        992 => "11111111",
        993 => "00010100",
        994 => "00010100",
        995 => "00010100",
        996 => "00010100",
        997 => "00010100",
        998 => "00010100",
        999 => "00010100",
        1000 => "00010100",
        1001 => "00010100",
        1002 => "00010100",
        1003 => "00010100",
        1004 => "00010100",
        1005 => "00010100",
        1006 => "00010100",
        1007 => "00010100",
        1008 => "00010100",
        1009 => "00010100",
        1010 => "00010100",
        1011 => "00010100",
        1012 => "00010100",
        1013 => "00010100",
        1014 => "00010100",
        1015 => "00010100",
        1016 => "00010100",
        1017 => "00010100",
        1018 => "00010100",
        1019 => "00010100",
        1020 => "00010100",
        1021 => "00010100",
        1022 => "00010100",
        1023 => "00010100",
        1024 => "00010100",
        1025 => "00010100",
        1026 => "00010100",
        1027 => "00010100",
        1028 => "00010100",
        1029 => "00010100",
        1030 => "00010100",
        1031 => "00010100",
        1032 => "00010100",
        1033 => "00010100",
        1034 => "00010100",
        1035 => "00010100",
        1036 => "00010100",
        1037 => "00010100",
        1038 => "00010100",
        1039 => "00010100",
        1040 => "00010100",
        1041 => "00010100",
        1042 => "00010100",
        1043 => "00010100",
        1044 => "00010100",
        1045 => "00000001",
        1046 => "00000001",
        1047 => "00000001",
        1048 => "00000001",
        1049 => "00000001",
        1050 => "00000001",
        1051 => "00000001",
        1052 => "00000001",
        1053 => "00000001",
        1054 => "00000001",
        1055 => "00000001",
        1056 => "00000001",
        1057 => "00000001",
        1058 => "00000001",
        1059 => "00000001",
        1060 => "00000001",
        1061 => "00000001",
        1062 => "00000001",
        1063 => "00000001",
        1064 => "00000001",
        1065 => "00000001",
        1066 => "00000001",
        1067 => "00000001",
        1068 => "00000001",
        1069 => "00000001",
        1070 => "00000001",
        1071 => "00000001",
        1072 => "00000001",
        1073 => "00000001",
        1074 => "00000001",
        1075 => "00000001",
        1076 => "00000001",
        1077 => "00000001",
        1078 => "00000001",
        1079 => "00000001",
        1080 => "00000001",
        1081 => "00000001",
        1082 => "00000001",
        1083 => "00000001",
        1084 => "00000001",
        1085 => "00000001",
        1086 => "00000001",
        1087 => "00000001",
        1088 => "00000001",
        1089 => "00000001",
        1090 => "00000001",
        1091 => "00000001",
        1092 => "00000001",
        1093 => "00000001",
        1094 => "00000001",
        1095 => "00000001",
        1096 => "00000001",
        1097 => "11111111",
        1098 => "11111111",
        1099 => "00000001",
        1100 => "00000001",
        1101 => "11111111",
        1102 => "11111111",
        1103 => "00010100",
        1104 => "00010100",
        1105 => "00010100",
        1106 => "00010100",
        1107 => "00010100",
        1108 => "00010100",
        1109 => "00010100",
        1110 => "00010100",
        1111 => "00010100",
        1112 => "00010100",
        1113 => "00010100",
        1114 => "00010100",
        1115 => "00010100",
        1116 => "00010101",
        1117 => "11011111",
        1118 => "11011101",
        1119 => "00010100",
        1120 => "00010100",
        1121 => "00010100",
        1122 => "00010100",
        1123 => "10011111",
        1124 => "11111111",
        1125 => "11111111",
        1126 => "11111111",
        1127 => "11111111",
        1128 => "11011001",
        1129 => "10111111",
        1130 => "11111101",
        1131 => "00010100",
        1132 => "00010100",
        1133 => "00010101",
        1134 => "11011111",
        1135 => "11011101",
        1136 => "01111111",
        1137 => "11111111",
        1138 => "11111111",
        1139 => "11111111",
        1140 => "11111111",
        1141 => "10111000",
        1142 => "00010100",
        1143 => "00010100",
        1144 => "00010100",
        1145 => "00010100",
        1146 => "00010100",
        1147 => "00010100",
        1148 => "00010100",
        1149 => "00010100",
        1150 => "00010100",
        1151 => "00010100",
        1152 => "00010100",
        1153 => "00010100",
        1154 => "00010100",
        1155 => "00000001",
        1156 => "00000001",
        1157 => "00000001",
        1158 => "00000001",
        1159 => "00000001",
        1160 => "00000001",
        1161 => "00000001",
        1162 => "00000001",
        1163 => "00000001",
        1164 => "00000001",
        1165 => "00000001",
        1166 => "00000001",
        1167 => "00000001",
        1168 => "00000001",
        1169 => "00000001",
        1170 => "00000001",
        1171 => "00000001",
        1172 => "00010011",
        1173 => "11111111",
        1174 => "11111111",
        1175 => "11111111",
        1176 => "10101101",
        1177 => "00000001",
        1178 => "00001110",
        1179 => "11011111",
        1180 => "11111111",
        1181 => "11111111",
        1182 => "11111111",
        1183 => "11010110",
        1184 => "00000001",
        1185 => "10011011",
        1186 => "11111111",
        1187 => "11111111",
        1188 => "11111111",
        1189 => "11111111",
        1190 => "10000001",
        1191 => "00000001",
        1192 => "00000001",
        1193 => "00000001",
        1194 => "00000001",
        1195 => "00000001",
        1196 => "00000001",
        1197 => "00000001",
        1198 => "00000001",
        1199 => "00000001",
        1200 => "00000001",
        1201 => "00000001",
        1202 => "00000001",
        1203 => "00000001",
        1204 => "00000001",
        1205 => "00000001",
        1206 => "00000001",
        1207 => "11111111",
        1208 => "11111111",
        1209 => "00000001",
        1210 => "00000001",
        1211 => "11111111",
        1212 => "11111111",
        1213 => "00010100",
        1214 => "00010100",
        1215 => "00010100",
        1216 => "00010100",
        1217 => "00010100",
        1218 => "00010100",
        1219 => "00010100",
        1220 => "00010100",
        1221 => "00010100",
        1222 => "00010100",
        1223 => "00010100",
        1224 => "00010100",
        1225 => "00010100",
        1226 => "00010101",
        1227 => "11011111",
        1228 => "11011101",
        1229 => "00010100",
        1230 => "00010100",
        1231 => "00010100",
        1232 => "00010100",
        1233 => "00010100",
        1234 => "00010101",
        1235 => "11011111",
        1236 => "11011101",
        1237 => "00010100",
        1238 => "00010100",
        1239 => "10011111",
        1240 => "11111110",
        1241 => "10010100",
        1242 => "00010100",
        1243 => "00011010",
        1244 => "11111111",
        1245 => "10111000",
        1246 => "01111111",
        1247 => "11111110",
        1248 => "10010100",
        1249 => "00010100",
        1250 => "00010100",
        1251 => "00010100",
        1252 => "00010100",
        1253 => "00010100",
        1254 => "00010100",
        1255 => "00010100",
        1256 => "00010100",
        1257 => "00010100",
        1258 => "00010100",
        1259 => "00010100",
        1260 => "00010100",
        1261 => "00010100",
        1262 => "00010100",
        1263 => "00010100",
        1264 => "00010100",
        1265 => "00000001",
        1266 => "00000001",
        1267 => "00000001",
        1268 => "00000001",
        1269 => "00000001",
        1270 => "00000001",
        1271 => "00000001",
        1272 => "00000001",
        1273 => "00000001",
        1274 => "00000001",
        1275 => "00000001",
        1276 => "00000001",
        1277 => "00000001",
        1278 => "00000001",
        1279 => "00000001",
        1280 => "00000001",
        1281 => "00001110",
        1282 => "11011111",
        1283 => "11010001",
        1284 => "00000001",
        1285 => "10011011",
        1286 => "11111010",
        1287 => "01100001",
        1288 => "00001110",
        1289 => "11011111",
        1290 => "11010001",
        1291 => "00000001",
        1292 => "00000001",
        1293 => "00000001",
        1294 => "00000001",
        1295 => "10011011",
        1296 => "11111010",
        1297 => "01100001",
        1298 => "00000001",
        1299 => "00000001",
        1300 => "00000001",
        1301 => "00000001",
        1302 => "00000001",
        1303 => "00000001",
        1304 => "00000001",
        1305 => "00000001",
        1306 => "00000001",
        1307 => "00000001",
        1308 => "00000001",
        1309 => "00000001",
        1310 => "00000001",
        1311 => "00000001",
        1312 => "00000001",
        1313 => "00000001",
        1314 => "00000001",
        1315 => "00000001",
        1316 => "00000001",
        1317 => "11111111",
        1318 => "11111111",
        1319 => "00000001",
        1320 => "00000001",
        1321 => "11111111",
        1322 => "11111111",
        1323 => "00010100",
        1324 => "00010100",
        1325 => "00010100",
        1326 => "00010100",
        1327 => "00010100",
        1328 => "00010100",
        1329 => "00010100",
        1330 => "00010100",
        1331 => "00010100",
        1332 => "00010100",
        1333 => "00010100",
        1334 => "00010100",
        1335 => "00010100",
        1336 => "00010101",
        1337 => "11011111",
        1338 => "11011101",
        1339 => "00010100",
        1340 => "00010100",
        1341 => "00010100",
        1342 => "00010100",
        1343 => "00010100",
        1344 => "00010101",
        1345 => "11011111",
        1346 => "11011101",
        1347 => "00010100",
        1348 => "00010100",
        1349 => "00011010",
        1350 => "11111111",
        1351 => "11011000",
        1352 => "00010100",
        1353 => "10011111",
        1354 => "11111110",
        1355 => "01110100",
        1356 => "01111111",
        1357 => "11111110",
        1358 => "10010100",
        1359 => "00010100",
        1360 => "00010100",
        1361 => "00010100",
        1362 => "00010100",
        1363 => "00010100",
        1364 => "00010100",
        1365 => "00010100",
        1366 => "00010100",
        1367 => "00010100",
        1368 => "00010100",
        1369 => "00010100",
        1370 => "00010100",
        1371 => "00010100",
        1372 => "00010100",
        1373 => "00010100",
        1374 => "00010100",
        1375 => "00000001",
        1376 => "00000001",
        1377 => "00000001",
        1378 => "00000001",
        1379 => "00000001",
        1380 => "00000001",
        1381 => "00000001",
        1382 => "00000001",
        1383 => "00000001",
        1384 => "00000001",
        1385 => "00000001",
        1386 => "00000001",
        1387 => "00000001",
        1388 => "00000001",
        1389 => "00000001",
        1390 => "00000001",
        1391 => "10011011",
        1392 => "11111010",
        1393 => "01100001",
        1394 => "00000001",
        1395 => "00010011",
        1396 => "11111111",
        1397 => "10101101",
        1398 => "00001110",
        1399 => "11011111",
        1400 => "11010001",
        1401 => "00000001",
        1402 => "00000001",
        1403 => "00000001",
        1404 => "00000001",
        1405 => "10011011",
        1406 => "11111010",
        1407 => "01100001",
        1408 => "00000001",
        1409 => "00000001",
        1410 => "00000001",
        1411 => "00000001",
        1412 => "00000001",
        1413 => "00000001",
        1414 => "00000001",
        1415 => "00000001",
        1416 => "00000001",
        1417 => "00000001",
        1418 => "00000001",
        1419 => "00000001",
        1420 => "00000001",
        1421 => "00000001",
        1422 => "00000001",
        1423 => "00000001",
        1424 => "00000001",
        1425 => "00000001",
        1426 => "00000001",
        1427 => "11111111",
        1428 => "11111111",
        1429 => "00000001",
        1430 => "00000001",
        1431 => "11111111",
        1432 => "11111111",
        1433 => "00010100",
        1434 => "00010100",
        1435 => "00010100",
        1436 => "00010100",
        1437 => "00010100",
        1438 => "00010100",
        1439 => "00010100",
        1440 => "00010100",
        1441 => "00010100",
        1442 => "00010100",
        1443 => "00010100",
        1444 => "00010100",
        1445 => "00010100",
        1446 => "00010101",
        1447 => "11011111",
        1448 => "11011101",
        1449 => "00010100",
        1450 => "00010100",
        1451 => "00010100",
        1452 => "00010100",
        1453 => "00010100",
        1454 => "00010101",
        1455 => "11011111",
        1456 => "11011101",
        1457 => "00010100",
        1458 => "00010100",
        1459 => "00010101",
        1460 => "11011111",
        1461 => "11011101",
        1462 => "00010101",
        1463 => "10111111",
        1464 => "11011101",
        1465 => "00010100",
        1466 => "01111111",
        1467 => "11111111",
        1468 => "11111111",
        1469 => "11111111",
        1470 => "11111110",
        1471 => "10010100",
        1472 => "00010100",
        1473 => "00010100",
        1474 => "00010100",
        1475 => "00010100",
        1476 => "00010100",
        1477 => "00010100",
        1478 => "00010100",
        1479 => "00010100",
        1480 => "00010100",
        1481 => "00010100",
        1482 => "00010100",
        1483 => "00010100",
        1484 => "00010100",
        1485 => "00000001",
        1486 => "00000001",
        1487 => "00000001",
        1488 => "00000001",
        1489 => "00000001",
        1490 => "00000001",
        1491 => "00000001",
        1492 => "00000001",
        1493 => "00000001",
        1494 => "00000001",
        1495 => "00000001",
        1496 => "00000001",
        1497 => "00000001",
        1498 => "00000001",
        1499 => "00000001",
        1500 => "00000001",
        1501 => "10011011",
        1502 => "11111010",
        1503 => "01100001",
        1504 => "00000001",
        1505 => "00001110",
        1506 => "11011111",
        1507 => "11010001",
        1508 => "00001110",
        1509 => "11011111",
        1510 => "11010001",
        1511 => "00000001",
        1512 => "00000001",
        1513 => "00000001",
        1514 => "00000001",
        1515 => "10011011",
        1516 => "11111010",
        1517 => "01100001",
        1518 => "00000001",
        1519 => "00000001",
        1520 => "00000001",
        1521 => "00000001",
        1522 => "00000001",
        1523 => "00000001",
        1524 => "00000001",
        1525 => "00000001",
        1526 => "00000001",
        1527 => "00000001",
        1528 => "00000001",
        1529 => "00000001",
        1530 => "00000001",
        1531 => "00000001",
        1532 => "00000001",
        1533 => "00000001",
        1534 => "00000001",
        1535 => "00000001",
        1536 => "00000001",
        1537 => "11111111",
        1538 => "11111111",
        1539 => "00000001",
        1540 => "00000001",
        1541 => "11111111",
        1542 => "11111111",
        1543 => "00010100",
        1544 => "00010100",
        1545 => "00010100",
        1546 => "00010100",
        1547 => "00010100",
        1548 => "00010100",
        1549 => "00010100",
        1550 => "00010100",
        1551 => "00010100",
        1552 => "00010100",
        1553 => "00010100",
        1554 => "00010100",
        1555 => "00010100",
        1556 => "00010101",
        1557 => "11011111",
        1558 => "11011101",
        1559 => "00010100",
        1560 => "00010100",
        1561 => "00010100",
        1562 => "00010100",
        1563 => "00010100",
        1564 => "00010101",
        1565 => "11011111",
        1566 => "11011101",
        1567 => "00010100",
        1568 => "00010100",
        1569 => "00010100",
        1570 => "10011111",
        1571 => "11111110",
        1572 => "01111010",
        1573 => "11011111",
        1574 => "11011000",
        1575 => "00010100",
        1576 => "01111111",
        1577 => "11111110",
        1578 => "10010100",
        1579 => "00010100",
        1580 => "00010100",
        1581 => "00010100",
        1582 => "00010100",
        1583 => "00010100",
        1584 => "00010100",
        1585 => "00010100",
        1586 => "00010100",
        1587 => "00010100",
        1588 => "00010100",
        1589 => "00010100",
        1590 => "00010100",
        1591 => "00010100",
        1592 => "00010100",
        1593 => "00010100",
        1594 => "00010100",
        1595 => "00000001",
        1596 => "00000001",
        1597 => "00000001",
        1598 => "00000001",
        1599 => "00000001",
        1600 => "00000001",
        1601 => "00000001",
        1602 => "00000001",
        1603 => "00000001",
        1604 => "00000001",
        1605 => "00000001",
        1606 => "00000001",
        1607 => "00000001",
        1608 => "00000001",
        1609 => "00000001",
        1610 => "00000001",
        1611 => "10011011",
        1612 => "11111010",
        1613 => "01100001",
        1614 => "00000001",
        1615 => "00001110",
        1616 => "11011111",
        1617 => "11010001",
        1618 => "00001110",
        1619 => "11011111",
        1620 => "11111111",
        1621 => "11111111",
        1622 => "11111111",
        1623 => "11010001",
        1624 => "00000001",
        1625 => "10011011",
        1626 => "11111111",
        1627 => "11111111",
        1628 => "11111111",
        1629 => "11111010",
        1630 => "01100001",
        1631 => "00000001",
        1632 => "00000001",
        1633 => "00000001",
        1634 => "00000001",
        1635 => "00000001",
        1636 => "00000001",
        1637 => "00000001",
        1638 => "00000001",
        1639 => "00000001",
        1640 => "00000001",
        1641 => "00000001",
        1642 => "00000001",
        1643 => "00000001",
        1644 => "00000001",
        1645 => "00000001",
        1646 => "00000001",
        1647 => "11111111",
        1648 => "11111111",
        1649 => "00000001",
        1650 => "00000001",
        1651 => "11111111",
        1652 => "11111111",
        1653 => "00010100",
        1654 => "00010100",
        1655 => "00010100",
        1656 => "00010100",
        1657 => "00010100",
        1658 => "00010100",
        1659 => "00010100",
        1660 => "00010100",
        1661 => "00010100",
        1662 => "00010100",
        1663 => "00010100",
        1664 => "00010100",
        1665 => "00010100",
        1666 => "00010101",
        1667 => "11011111",
        1668 => "11011101",
        1669 => "00010100",
        1670 => "00010100",
        1671 => "00010100",
        1672 => "00010100",
        1673 => "00010100",
        1674 => "00010101",
        1675 => "11011111",
        1676 => "11011101",
        1677 => "00010100",
        1678 => "00010100",
        1679 => "00010100",
        1680 => "00011010",
        1681 => "11111111",
        1682 => "11011111",
        1683 => "11111110",
        1684 => "10010100",
        1685 => "00010100",
        1686 => "01111111",
        1687 => "11111110",
        1688 => "10010100",
        1689 => "00010100",
        1690 => "00010100",
        1691 => "00010100",
        1692 => "00010100",
        1693 => "00010100",
        1694 => "00010100",
        1695 => "00010100",
        1696 => "00010100",
        1697 => "00010100",
        1698 => "00010100",
        1699 => "00010100",
        1700 => "00010100",
        1701 => "00010100",
        1702 => "00010100",
        1703 => "00010100",
        1704 => "00010100",
        1705 => "00000001",
        1706 => "00000001",
        1707 => "00000001",
        1708 => "00000001",
        1709 => "00000001",
        1710 => "00000001",
        1711 => "00000001",
        1712 => "00000001",
        1713 => "00000001",
        1714 => "00000001",
        1715 => "00000001",
        1716 => "00000001",
        1717 => "00000001",
        1718 => "00000001",
        1719 => "00000001",
        1720 => "00000001",
        1721 => "10011011",
        1722 => "11111010",
        1723 => "01100001",
        1724 => "00000001",
        1725 => "00001110",
        1726 => "11011111",
        1727 => "10101101",
        1728 => "00001110",
        1729 => "11011111",
        1730 => "11010001",
        1731 => "00000001",
        1732 => "00000001",
        1733 => "00000001",
        1734 => "00000001",
        1735 => "10011011",
        1736 => "11111010",
        1737 => "01100001",
        1738 => "00000001",
        1739 => "00000001",
        1740 => "00000001",
        1741 => "00000001",
        1742 => "00000001",
        1743 => "00000001",
        1744 => "00000001",
        1745 => "00000001",
        1746 => "00000001",
        1747 => "00000001",
        1748 => "00000001",
        1749 => "00000001",
        1750 => "00000001",
        1751 => "00000001",
        1752 => "00000001",
        1753 => "00000001",
        1754 => "00000001",
        1755 => "00000001",
        1756 => "00000001",
        1757 => "11111111",
        1758 => "11111111",
        1759 => "00000001",
        1760 => "00000001",
        1761 => "11111111",
        1762 => "11111111",
        1763 => "00010100",
        1764 => "00010100",
        1765 => "00010100",
        1766 => "00010100",
        1767 => "00010100",
        1768 => "00010100",
        1769 => "00010100",
        1770 => "00010100",
        1771 => "00010100",
        1772 => "00010100",
        1773 => "00010100",
        1774 => "00010100",
        1775 => "00010100",
        1776 => "00010101",
        1777 => "11011111",
        1778 => "11011101",
        1779 => "00010100",
        1780 => "00010100",
        1781 => "00010100",
        1782 => "00010100",
        1783 => "00010100",
        1784 => "00010101",
        1785 => "11011111",
        1786 => "11011101",
        1787 => "00010100",
        1788 => "00010100",
        1789 => "00010100",
        1790 => "00011010",
        1791 => "11011111",
        1792 => "11111111",
        1793 => "11111101",
        1794 => "00010100",
        1795 => "00010100",
        1796 => "01111111",
        1797 => "11111110",
        1798 => "10010100",
        1799 => "00010100",
        1800 => "00010100",
        1801 => "00010100",
        1802 => "00010100",
        1803 => "00010100",
        1804 => "00010100",
        1805 => "00010100",
        1806 => "00010100",
        1807 => "00010100",
        1808 => "00010100",
        1809 => "00010100",
        1810 => "00010100",
        1811 => "00010100",
        1812 => "00010100",
        1813 => "00010100",
        1814 => "00010100",
        1815 => "00000001",
        1816 => "00000001",
        1817 => "00000001",
        1818 => "00000001",
        1819 => "00000001",
        1820 => "00000001",
        1821 => "00000001",
        1822 => "00000001",
        1823 => "00000001",
        1824 => "00000001",
        1825 => "00000001",
        1826 => "00000001",
        1827 => "00000001",
        1828 => "00000001",
        1829 => "00000001",
        1830 => "00000001",
        1831 => "00010011",
        1832 => "11111111",
        1833 => "11010001",
        1834 => "00000001",
        1835 => "10011011",
        1836 => "11111010",
        1837 => "01100001",
        1838 => "00001110",
        1839 => "11011111",
        1840 => "11010001",
        1841 => "00000001",
        1842 => "00000001",
        1843 => "00000001",
        1844 => "00000001",
        1845 => "10011011",
        1846 => "11111010",
        1847 => "01100001",
        1848 => "00000001",
        1849 => "00000001",
        1850 => "00000001",
        1851 => "00000001",
        1852 => "00000001",
        1853 => "00000001",
        1854 => "00000001",
        1855 => "00000001",
        1856 => "00000001",
        1857 => "00000001",
        1858 => "00000001",
        1859 => "00000001",
        1860 => "00000001",
        1861 => "00000001",
        1862 => "00000001",
        1863 => "00000001",
        1864 => "00000001",
        1865 => "00000001",
        1866 => "00000001",
        1867 => "11111111",
        1868 => "11111111",
        1869 => "00000001",
        1870 => "00000001",
        1871 => "11111111",
        1872 => "11111111",
        1873 => "00010100",
        1874 => "00010100",
        1875 => "00010100",
        1876 => "00010100",
        1877 => "00010100",
        1878 => "00010100",
        1879 => "00010100",
        1880 => "00010100",
        1881 => "00010100",
        1882 => "00010100",
        1883 => "00010100",
        1884 => "00010100",
        1885 => "00010100",
        1886 => "00010101",
        1887 => "11011111",
        1888 => "11111111",
        1889 => "11111111",
        1890 => "11111111",
        1891 => "11111101",
        1892 => "00010100",
        1893 => "10011111",
        1894 => "11111111",
        1895 => "11111111",
        1896 => "11111111",
        1897 => "11111111",
        1898 => "11011000",
        1899 => "00010100",
        1900 => "00010101",
        1901 => "10111111",
        1902 => "11111111",
        1903 => "11011000",
        1904 => "00010100",
        1905 => "00010100",
        1906 => "01111111",
        1907 => "11111111",
        1908 => "11111111",
        1909 => "11111111",
        1910 => "11111111",
        1911 => "10111000",
        1912 => "00010100",
        1913 => "00010100",
        1914 => "00010100",
        1915 => "00010100",
        1916 => "00010100",
        1917 => "00010100",
        1918 => "00010100",
        1919 => "00010100",
        1920 => "00010100",
        1921 => "00010100",
        1922 => "00010100",
        1923 => "00010100",
        1924 => "00010100",
        1925 => "00000001",
        1926 => "00000001",
        1927 => "00000001",
        1928 => "00000001",
        1929 => "00000001",
        1930 => "00000001",
        1931 => "00000001",
        1932 => "00000001",
        1933 => "00000001",
        1934 => "00000001",
        1935 => "00000001",
        1936 => "00000001",
        1937 => "00000001",
        1938 => "00000001",
        1939 => "00000001",
        1940 => "00000001",
        1941 => "00000001",
        1942 => "01110111",
        1943 => "11111111",
        1944 => "11111111",
        1945 => "11111111",
        1946 => "10000001",
        1947 => "00000001",
        1948 => "00001110",
        1949 => "11011111",
        1950 => "11010001",
        1951 => "00000001",
        1952 => "00000001",
        1953 => "00000001",
        1954 => "00000001",
        1955 => "10011011",
        1956 => "11111010",
        1957 => "01100001",
        1958 => "00000001",
        1959 => "00000001",
        1960 => "00000001",
        1961 => "00000001",
        1962 => "00000001",
        1963 => "00000001",
        1964 => "00000001",
        1965 => "00000001",
        1966 => "00000001",
        1967 => "00000001",
        1968 => "00000001",
        1969 => "00000001",
        1970 => "00000001",
        1971 => "00000001",
        1972 => "00000001",
        1973 => "00000001",
        1974 => "00000001",
        1975 => "00000001",
        1976 => "00000001",
        1977 => "11111111",
        1978 => "11111111",
        1979 => "00000001",
        1980 => "00000001",
        1981 => "11111111",
        1982 => "11111111",
        1983 => "00010100",
        1984 => "00010100",
        1985 => "00010100",
        1986 => "00010100",
        1987 => "00010100",
        1988 => "00010100",
        1989 => "00010100",
        1990 => "00010100",
        1991 => "00010100",
        1992 => "00010100",
        1993 => "00010100",
        1994 => "00010100",
        1995 => "00010100",
        1996 => "00010100",
        1997 => "00010100",
        1998 => "00010100",
        1999 => "00010100",
        2000 => "00010100",
        2001 => "00010100",
        2002 => "00010100",
        2003 => "00010100",
        2004 => "00010100",
        2005 => "00010100",
        2006 => "00010100",
        2007 => "00010100",
        2008 => "00010100",
        2009 => "00010100",
        2010 => "00010100",
        2011 => "00010100",
        2012 => "00010100",
        2013 => "00010100",
        2014 => "00010100",
        2015 => "00010100",
        2016 => "00010100",
        2017 => "00010100",
        2018 => "00010100",
        2019 => "00010100",
        2020 => "00010100",
        2021 => "00010100",
        2022 => "00010100",
        2023 => "00010100",
        2024 => "00010100",
        2025 => "00010100",
        2026 => "00010100",
        2027 => "00010100",
        2028 => "00010100",
        2029 => "00010100",
        2030 => "00010100",
        2031 => "00010100",
        2032 => "00010100",
        2033 => "00010100",
        2034 => "00010100",
        2035 => "00000001",
        2036 => "00000001",
        2037 => "00000001",
        2038 => "00000001",
        2039 => "00000001",
        2040 => "00000001",
        2041 => "00000001",
        2042 => "00000001",
        2043 => "00000001",
        2044 => "00000001",
        2045 => "00000001",
        2046 => "00000001",
        2047 => "00000001",
        2048 => "00000001",
        2049 => "00000001",
        2050 => "00000001",
        2051 => "00000001",
        2052 => "00000001",
        2053 => "00000001",
        2054 => "00000001",
        2055 => "00000001",
        2056 => "00000001",
        2057 => "00000001",
        2058 => "00000001",
        2059 => "00000001",
        2060 => "00000001",
        2061 => "00000001",
        2062 => "00000001",
        2063 => "00000001",
        2064 => "00000001",
        2065 => "00000001",
        2066 => "00000001",
        2067 => "00000001",
        2068 => "00000001",
        2069 => "00000001",
        2070 => "00000001",
        2071 => "00000001",
        2072 => "00000001",
        2073 => "00000001",
        2074 => "00000001",
        2075 => "00000001",
        2076 => "00000001",
        2077 => "00000001",
        2078 => "00000001",
        2079 => "00000001",
        2080 => "00000001",
        2081 => "00000001",
        2082 => "00000001",
        2083 => "00000001",
        2084 => "00000001",
        2085 => "00000001",
        2086 => "00000001",
        2087 => "11111111",
        2088 => "11111111",
        2089 => "00000001",
        2090 => "00000001",
        2091 => "11111111",
        2092 => "11111111",
        2093 => "00010100",
        2094 => "00010100",
        2095 => "00010100",
        2096 => "00010100",
        2097 => "00010100",
        2098 => "00010100",
        2099 => "00010100",
        2100 => "00010100",
        2101 => "00010100",
        2102 => "00010100",
        2103 => "00010100",
        2104 => "00010100",
        2105 => "00010100",
        2106 => "00010100",
        2107 => "00010100",
        2108 => "00010100",
        2109 => "00010100",
        2110 => "00010100",
        2111 => "00010100",
        2112 => "00010100",
        2113 => "00010100",
        2114 => "00010100",
        2115 => "00010100",
        2116 => "00010100",
        2117 => "00010100",
        2118 => "00010100",
        2119 => "00010100",
        2120 => "00010100",
        2121 => "00010100",
        2122 => "00010100",
        2123 => "00010100",
        2124 => "00010100",
        2125 => "00010100",
        2126 => "00010100",
        2127 => "00010100",
        2128 => "00010100",
        2129 => "00010100",
        2130 => "00010100",
        2131 => "00010100",
        2132 => "00010100",
        2133 => "00010100",
        2134 => "00010100",
        2135 => "00010100",
        2136 => "00010100",
        2137 => "00010100",
        2138 => "00010100",
        2139 => "00010100",
        2140 => "00010100",
        2141 => "00010100",
        2142 => "00010100",
        2143 => "00010100",
        2144 => "00010100",
        2145 => "00000001",
        2146 => "00000001",
        2147 => "00000001",
        2148 => "00000001",
        2149 => "00000001",
        2150 => "00000001",
        2151 => "00000001",
        2152 => "00000001",
        2153 => "00000001",
        2154 => "00000001",
        2155 => "00000001",
        2156 => "00000001",
        2157 => "00000001",
        2158 => "00000001",
        2159 => "00000001",
        2160 => "00000001",
        2161 => "00000001",
        2162 => "00000001",
        2163 => "00000001",
        2164 => "00000001",
        2165 => "00000001",
        2166 => "00000001",
        2167 => "00000001",
        2168 => "00000001",
        2169 => "00000001",
        2170 => "00000001",
        2171 => "00000001",
        2172 => "00000001",
        2173 => "00000001",
        2174 => "00000001",
        2175 => "00000001",
        2176 => "00000001",
        2177 => "00000001",
        2178 => "00000001",
        2179 => "00000001",
        2180 => "00000001",
        2181 => "00000001",
        2182 => "00000001",
        2183 => "00000001",
        2184 => "00000001",
        2185 => "00000001",
        2186 => "00000001",
        2187 => "00000001",
        2188 => "00000001",
        2189 => "00000001",
        2190 => "00000001",
        2191 => "00000001",
        2192 => "00000001",
        2193 => "00000001",
        2194 => "00000001",
        2195 => "00000001",
        2196 => "00000001",
        2197 => "11111111",
        2198 => "11111111",
        2199 => "00000001",
        2200 => "00000001",
        2201 => "11111111",
        2202 => "11111111",
        2203 => "00010100",
        2204 => "00010100",
        2205 => "00010100",
        2206 => "00010100",
        2207 => "00010100",
        2208 => "00010100",
        2209 => "00010100",
        2210 => "00010100",
        2211 => "00010100",
        2212 => "00010100",
        2213 => "00010100",
        2214 => "00010100",
        2215 => "00010100",
        2216 => "00010100",
        2217 => "00010100",
        2218 => "00010100",
        2219 => "00010100",
        2220 => "00010100",
        2221 => "00010100",
        2222 => "00010100",
        2223 => "00010100",
        2224 => "00010100",
        2225 => "00010100",
        2226 => "00010100",
        2227 => "00010100",
        2228 => "00010100",
        2229 => "00010100",
        2230 => "00010100",
        2231 => "00010100",
        2232 => "00010100",
        2233 => "00010100",
        2234 => "00010100",
        2235 => "00010100",
        2236 => "00010100",
        2237 => "00010100",
        2238 => "00010100",
        2239 => "00010100",
        2240 => "00010100",
        2241 => "00010100",
        2242 => "00010100",
        2243 => "00010100",
        2244 => "00010100",
        2245 => "00010100",
        2246 => "00010100",
        2247 => "00010100",
        2248 => "00010100",
        2249 => "00010100",
        2250 => "00010100",
        2251 => "00010100",
        2252 => "00010100",
        2253 => "00010100",
        2254 => "00010100",
        2255 => "00000001",
        2256 => "00000001",
        2257 => "00000001",
        2258 => "00000001",
        2259 => "00000001",
        2260 => "00000001",
        2261 => "00000001",
        2262 => "00000001",
        2263 => "00000001",
        2264 => "00000001",
        2265 => "00000001",
        2266 => "00000001",
        2267 => "00000001",
        2268 => "00000001",
        2269 => "00000001",
        2270 => "00000001",
        2271 => "00000001",
        2272 => "00000001",
        2273 => "00000001",
        2274 => "00000001",
        2275 => "00000001",
        2276 => "00000001",
        2277 => "00000001",
        2278 => "00000001",
        2279 => "00000001",
        2280 => "00000001",
        2281 => "00000001",
        2282 => "00000001",
        2283 => "00000001",
        2284 => "00000001",
        2285 => "00000001",
        2286 => "00000001",
        2287 => "00000001",
        2288 => "00000001",
        2289 => "00000001",
        2290 => "00000001",
        2291 => "00000001",
        2292 => "00000001",
        2293 => "00000001",
        2294 => "00000001",
        2295 => "00000001",
        2296 => "00000001",
        2297 => "00000001",
        2298 => "00000001",
        2299 => "00000001",
        2300 => "00000001",
        2301 => "00000001",
        2302 => "00000001",
        2303 => "00000001",
        2304 => "00000001",
        2305 => "00000001",
        2306 => "00000001",
        2307 => "11111111",
        2308 => "11111111",
        2309 => "00000001",
        2310 => "00000001",
        2311 => "11111111",
        2312 => "11111111",
        2313 => "00010100",
        2314 => "00010100",
        2315 => "00010100",
        2316 => "00010100",
        2317 => "00010100",
        2318 => "00010100",
        2319 => "00010100",
        2320 => "00010100",
        2321 => "00010100",
        2322 => "00010100",
        2323 => "00010100",
        2324 => "00010100",
        2325 => "00010100",
        2326 => "00010100",
        2327 => "00010100",
        2328 => "00010100",
        2329 => "00010100",
        2330 => "00010100",
        2331 => "00010100",
        2332 => "00010100",
        2333 => "00010100",
        2334 => "00010100",
        2335 => "00010100",
        2336 => "00010100",
        2337 => "00010100",
        2338 => "00010100",
        2339 => "00010100",
        2340 => "00010100",
        2341 => "00010100",
        2342 => "00010100",
        2343 => "00010100",
        2344 => "00010100",
        2345 => "00010100",
        2346 => "00010100",
        2347 => "00010100",
        2348 => "00010100",
        2349 => "00010100",
        2350 => "00010100",
        2351 => "00010100",
        2352 => "00010100",
        2353 => "00010100",
        2354 => "00010100",
        2355 => "00010100",
        2356 => "00010100",
        2357 => "00010100",
        2358 => "00010100",
        2359 => "00010100",
        2360 => "00010100",
        2361 => "00010100",
        2362 => "00010100",
        2363 => "00010100",
        2364 => "00010100",
        2365 => "00000001",
        2366 => "00000001",
        2367 => "00000001",
        2368 => "00000001",
        2369 => "00000001",
        2370 => "00000001",
        2371 => "00000001",
        2372 => "00000001",
        2373 => "00000001",
        2374 => "00000001",
        2375 => "00000001",
        2376 => "00000001",
        2377 => "00000001",
        2378 => "00000001",
        2379 => "00000001",
        2380 => "00000001",
        2381 => "00000001",
        2382 => "00000001",
        2383 => "00000001",
        2384 => "00000001",
        2385 => "00000001",
        2386 => "00000001",
        2387 => "00000001",
        2388 => "00000001",
        2389 => "00000001",
        2390 => "00000001",
        2391 => "00000001",
        2392 => "00000001",
        2393 => "00000001",
        2394 => "00000001",
        2395 => "00000001",
        2396 => "00000001",
        2397 => "00000001",
        2398 => "00000001",
        2399 => "00000001",
        2400 => "00000001",
        2401 => "00000001",
        2402 => "00000001",
        2403 => "00000001",
        2404 => "00000001",
        2405 => "00000001",
        2406 => "00000001",
        2407 => "00000001",
        2408 => "00000001",
        2409 => "00000001",
        2410 => "00000001",
        2411 => "00000001",
        2412 => "00000001",
        2413 => "00000001",
        2414 => "00000001",
        2415 => "00000001",
        2416 => "00000001",
        2417 => "11111111",
        2418 => "11111111",
        2419 => "00000001",
        2420 => "00000001",
        2421 => "11111111",
        2422 => "11111111",
        2423 => "00010100",
        2424 => "00010100",
        2425 => "00010100",
        2426 => "00010100",
        2427 => "00010100",
        2428 => "00010100",
        2429 => "00010100",
        2430 => "00010100",
        2431 => "00010100",
        2432 => "00010100",
        2433 => "00010100",
        2434 => "00010100",
        2435 => "00010100",
        2436 => "00010100",
        2437 => "00010100",
        2438 => "00010100",
        2439 => "00010100",
        2440 => "00010100",
        2441 => "00010100",
        2442 => "00010100",
        2443 => "00010100",
        2444 => "00010100",
        2445 => "00010100",
        2446 => "00010100",
        2447 => "00010100",
        2448 => "00010100",
        2449 => "00010100",
        2450 => "00010100",
        2451 => "00010100",
        2452 => "00010100",
        2453 => "00010100",
        2454 => "00010100",
        2455 => "00010100",
        2456 => "00010100",
        2457 => "00010100",
        2458 => "00010100",
        2459 => "00010100",
        2460 => "00010100",
        2461 => "00010100",
        2462 => "00010100",
        2463 => "00010100",
        2464 => "00010100",
        2465 => "00010100",
        2466 => "00010100",
        2467 => "00010100",
        2468 => "00010100",
        2469 => "00010100",
        2470 => "00010100",
        2471 => "00010100",
        2472 => "00010100",
        2473 => "00010100",
        2474 => "00010100",
        2475 => "00000001",
        2476 => "00000001",
        2477 => "00000001",
        2478 => "00000001",
        2479 => "00000001",
        2480 => "00000001",
        2481 => "00000001",
        2482 => "00000001",
        2483 => "00000001",
        2484 => "00000001",
        2485 => "00000001",
        2486 => "00000001",
        2487 => "00000001",
        2488 => "00000001",
        2489 => "00000001",
        2490 => "00000001",
        2491 => "00000001",
        2492 => "00000001",
        2493 => "00000001",
        2494 => "00000001",
        2495 => "00000001",
        2496 => "00000001",
        2497 => "00000001",
        2498 => "00000001",
        2499 => "00000001",
        2500 => "00000001",
        2501 => "00000001",
        2502 => "00000001",
        2503 => "00000001",
        2504 => "00000001",
        2505 => "00000001",
        2506 => "00000001",
        2507 => "00000001",
        2508 => "00000001",
        2509 => "00000001",
        2510 => "00000001",
        2511 => "00000001",
        2512 => "00000001",
        2513 => "00000001",
        2514 => "00000001",
        2515 => "00000001",
        2516 => "00000001",
        2517 => "00000001",
        2518 => "00000001",
        2519 => "00000001",
        2520 => "00000001",
        2521 => "00000001",
        2522 => "00000001",
        2523 => "00000001",
        2524 => "00000001",
        2525 => "00000001",
        2526 => "00000001",
        2527 => "11111111",
        2528 => "11111111",
        2529 => "00000001",
        2530 => "00000001",
        2531 => "11111111",
        2532 => "11111111",
        2533 => "00010100",
        2534 => "00010100",
        2535 => "00010100",
        2536 => "00010100",
        2537 => "00010100",
        2538 => "00010100",
        2539 => "00010100",
        2540 => "00010100",
        2541 => "00010100",
        2542 => "00010100",
        2543 => "00010100",
        2544 => "00010100",
        2545 => "00010100",
        2546 => "00010100",
        2547 => "00010100",
        2548 => "00010100",
        2549 => "00010100",
        2550 => "00010100",
        2551 => "00010100",
        2552 => "00010100",
        2553 => "00010100",
        2554 => "00010100",
        2555 => "00010100",
        2556 => "00010100",
        2557 => "00010100",
        2558 => "00010100",
        2559 => "00010100",
        2560 => "00010100",
        2561 => "00010100",
        2562 => "00010100",
        2563 => "00010100",
        2564 => "00010100",
        2565 => "00010100",
        2566 => "00010100",
        2567 => "00010100",
        2568 => "00010100",
        2569 => "00010100",
        2570 => "00010100",
        2571 => "00010100",
        2572 => "00010100",
        2573 => "00010100",
        2574 => "00010100",
        2575 => "00010100",
        2576 => "00010100",
        2577 => "00010100",
        2578 => "00010100",
        2579 => "00010100",
        2580 => "00010100",
        2581 => "00010100",
        2582 => "00010100",
        2583 => "00010100",
        2584 => "00010100",
        2585 => "00000001",
        2586 => "00000001",
        2587 => "00000001",
        2588 => "00000001",
        2589 => "00000001",
        2590 => "00000001",
        2591 => "00000001",
        2592 => "00000001",
        2593 => "00000001",
        2594 => "00000001",
        2595 => "00000001",
        2596 => "00000001",
        2597 => "00000001",
        2598 => "00000001",
        2599 => "00000001",
        2600 => "00000001",
        2601 => "00000001",
        2602 => "00000001",
        2603 => "00000001",
        2604 => "00000001",
        2605 => "00000001",
        2606 => "00000001",
        2607 => "00000001",
        2608 => "00000001",
        2609 => "00000001",
        2610 => "00000001",
        2611 => "00000001",
        2612 => "00000001",
        2613 => "00000001",
        2614 => "00000001",
        2615 => "00000001",
        2616 => "00000001",
        2617 => "00000001",
        2618 => "00000001",
        2619 => "00000001",
        2620 => "00000001",
        2621 => "00000001",
        2622 => "00000001",
        2623 => "00000001",
        2624 => "00000001",
        2625 => "00000001",
        2626 => "00000001",
        2627 => "00000001",
        2628 => "00000001",
        2629 => "00000001",
        2630 => "00000001",
        2631 => "00000001",
        2632 => "00000001",
        2633 => "00000001",
        2634 => "00000001",
        2635 => "00000001",
        2636 => "00000001",
        2637 => "11111111",
        2638 => "11111111",
        2639 => "00000001",
        2640 => "00000001",
        2641 => "10110110",
        2642 => "11111111",
        2643 => "01010001",
        2644 => "00010100",
        2645 => "00010100",
        2646 => "00010100",
        2647 => "00010100",
        2648 => "00010100",
        2649 => "00010100",
        2650 => "00010100",
        2651 => "00010100",
        2652 => "00010100",
        2653 => "00010100",
        2654 => "00010100",
        2655 => "00010100",
        2656 => "00010100",
        2657 => "00010100",
        2658 => "00010100",
        2659 => "00010100",
        2660 => "00010100",
        2661 => "00010100",
        2662 => "00010100",
        2663 => "00010100",
        2664 => "00010100",
        2665 => "00010100",
        2666 => "00010100",
        2667 => "00010100",
        2668 => "00010100",
        2669 => "00010100",
        2670 => "00010100",
        2671 => "00010100",
        2672 => "00010100",
        2673 => "00010100",
        2674 => "00010100",
        2675 => "00010100",
        2676 => "00010100",
        2677 => "00010100",
        2678 => "00010100",
        2679 => "00010100",
        2680 => "00010100",
        2681 => "00010100",
        2682 => "00010100",
        2683 => "00010100",
        2684 => "00010100",
        2685 => "00010100",
        2686 => "00010100",
        2687 => "00010100",
        2688 => "00010100",
        2689 => "00010100",
        2690 => "00010100",
        2691 => "00010100",
        2692 => "00010100",
        2693 => "00010100",
        2694 => "00010100",
        2695 => "00000001",
        2696 => "00000001",
        2697 => "00000001",
        2698 => "00000001",
        2699 => "00000001",
        2700 => "00000001",
        2701 => "00000001",
        2702 => "00000001",
        2703 => "00000001",
        2704 => "00000001",
        2705 => "00000001",
        2706 => "00000001",
        2707 => "00000001",
        2708 => "00000001",
        2709 => "00000001",
        2710 => "00000001",
        2711 => "00000001",
        2712 => "00000001",
        2713 => "00000001",
        2714 => "00000001",
        2715 => "00000001",
        2716 => "00000001",
        2717 => "00000001",
        2718 => "00000001",
        2719 => "00000001",
        2720 => "00000001",
        2721 => "00000001",
        2722 => "00000001",
        2723 => "00000001",
        2724 => "00000001",
        2725 => "00000001",
        2726 => "00000001",
        2727 => "00000001",
        2728 => "00000001",
        2729 => "00000001",
        2730 => "00000001",
        2731 => "00000001",
        2732 => "00000001",
        2733 => "00000001",
        2734 => "00000001",
        2735 => "00000001",
        2736 => "00000001",
        2737 => "00000001",
        2738 => "00000001",
        2739 => "00000001",
        2740 => "00000001",
        2741 => "00000001",
        2742 => "00000001",
        2743 => "00000001",
        2744 => "00000001",
        2745 => "00000001",
        2746 => "01001010",
        2747 => "11111111",
        2748 => "10110110",
        2749 => "00000001");
begin
    process(clk)
    begin
        if rising_edge(clk) then
            if rst = '1' then
                live <= (others => (others => '0'));
            else
                dout <= live(to_integer(unsigned(addr)));
            end if;
        end if;
    end process;


end Behavioral;

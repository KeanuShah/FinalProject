
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
entity View_Button is
    port(clk, rst: in std_logic;
         addr: in std_logic_vector(10 downto 0);
         dout: out std_logic_vector(7 downto 0));
    
end View_Button;

architecture Behavioral of View_Button is

    type mem is array (0 to 1733) of std_logic_vector(7 downto 0); 
    signal view: mem:= (
        0 => "00000001",
        1 => "00000001",
        2 => "00000001",
        3 => "00000000",
        4 => "00000001",
        5 => "00000001",
        6 => "00000000",
        7 => "00000000",
        8 => "00000000",
        9 => "00000000",
        10 => "00000000",
        11 => "00000000",
        12 => "00000000",
        13 => "00000000",
        14 => "00000000",
        15 => "00000000",
        16 => "00000000",
        17 => "00000000",
        18 => "00000000",
        19 => "00000000",
        20 => "00000000",
        21 => "00000000",
        22 => "00000000",
        23 => "00000000",
        24 => "00000000",
        25 => "00000000",
        26 => "00000000",
        27 => "00000000",
        28 => "00000000",
        29 => "00000000",
        30 => "00000000",
        31 => "00000000",
        32 => "00000000",
        33 => "00000000",
        34 => "00000000",
        35 => "00000000",
        36 => "00000000",
        37 => "00000000",
        38 => "00000000",
        39 => "00000000",
        40 => "00000001",
        41 => "00000001",
        42 => "00000000",
        43 => "00000000",
        44 => "00000000",
        45 => "00000000",
        46 => "00000001",
        47 => "00000001",
        48 => "00000000",
        49 => "00000001",
        50 => "00000001",
        51 => "00000001",
        52 => "00000001",
        53 => "00100101",
        54 => "10110111",
        55 => "11011111",
        56 => "11011111",
        57 => "11111111",
        58 => "11111111",
        59 => "11011111",
        60 => "11011111",
        61 => "11011111",
        62 => "11111111",
        63 => "11111111",
        64 => "11011111",
        65 => "11011111",
        66 => "11011111",
        67 => "11011111",
        68 => "11011111",
        69 => "11011111",
        70 => "11011111",
        71 => "11111111",
        72 => "11111111",
        73 => "11011111",
        74 => "11011111",
        75 => "11011111",
        76 => "11011111",
        77 => "11011111",
        78 => "11011111",
        79 => "11111111",
        80 => "11111111",
        81 => "11011111",
        82 => "11011111",
        83 => "11011111",
        84 => "11011111",
        85 => "11111111",
        86 => "11111111",
        87 => "11011111",
        88 => "11011111",
        89 => "11011111",
        90 => "11011111",
        91 => "11011111",
        92 => "11011111",
        93 => "11011111",
        94 => "11011111",
        95 => "11011111",
        96 => "11011111",
        97 => "11011011",
        98 => "10010011",
        99 => "00100101",
        100 => "00000000",
        101 => "00000001",
        102 => "00000001",
        103 => "00101001",
        104 => "11011111",
        105 => "11011111",
        106 => "10111111",
        107 => "10111111",
        108 => "11011110",
        109 => "10111110",
        110 => "10111110",
        111 => "10111110",
        112 => "10111110",
        113 => "10111110",
        114 => "10111110",
        115 => "10111110",
        116 => "10111110",
        117 => "10111110",
        118 => "10111110",
        119 => "10111110",
        120 => "10111110",
        121 => "10111110",
        122 => "10111110",
        123 => "11011110",
        124 => "10111110",
        125 => "10111110",
        126 => "10111110",
        127 => "10111110",
        128 => "10111111",
        129 => "10111111",
        130 => "10111110",
        131 => "10111110",
        132 => "10111110",
        133 => "10111110",
        134 => "10111110",
        135 => "10111110",
        136 => "10111110",
        137 => "10111110",
        138 => "10111110",
        139 => "10111110",
        140 => "10111110",
        141 => "10111111",
        142 => "10111111",
        143 => "10111111",
        144 => "10111110",
        145 => "10111110",
        146 => "10111110",
        147 => "11011110",
        148 => "11011111",
        149 => "11011111",
        150 => "10111011",
        151 => "00100101",
        152 => "00000001",
        153 => "00000000",
        154 => "10110111",
        155 => "11011111",
        156 => "10011001",
        157 => "00110000",
        158 => "00010000",
        159 => "00010000",
        160 => "00001100",
        161 => "00010000",
        162 => "00010000",
        163 => "00010000",
        164 => "00001100",
        165 => "00010000",
        166 => "00010000",
        167 => "00010000",
        168 => "00010000",
        169 => "00010000",
        170 => "00010000",
        171 => "00010000",
        172 => "00010000",
        173 => "00010000",
        174 => "00010000",
        175 => "00001100",
        176 => "00001100",
        177 => "00001100",
        178 => "00001100",
        179 => "00001100",
        180 => "00001100",
        181 => "00001100",
        182 => "00001100",
        183 => "00010000",
        184 => "00010000",
        185 => "00001100",
        186 => "00010000",
        187 => "00010000",
        188 => "00010000",
        189 => "00010000",
        190 => "00010000",
        191 => "00010000",
        192 => "00010000",
        193 => "00001100",
        194 => "00010000",
        195 => "00010000",
        196 => "00010000",
        197 => "00010000",
        198 => "00001100",
        199 => "00110000",
        200 => "10011010",
        201 => "11011111",
        202 => "10010011",
        203 => "00000001",
        204 => "00000101",
        205 => "11011111",
        206 => "10111111",
        207 => "00110000",
        208 => "00010000",
        209 => "00010000",
        210 => "00010000",
        211 => "00010000",
        212 => "00010000",
        213 => "00010000",
        214 => "00010000",
        215 => "00010000",
        216 => "00010000",
        217 => "00010000",
        218 => "00010000",
        219 => "00010000",
        220 => "00010000",
        221 => "00010000",
        222 => "00010000",
        223 => "00010000",
        224 => "00010000",
        225 => "00010000",
        226 => "00010000",
        227 => "00010000",
        228 => "00010000",
        229 => "00010000",
        230 => "00010000",
        231 => "00010000",
        232 => "00010000",
        233 => "00010000",
        234 => "00010000",
        235 => "00010000",
        236 => "00010000",
        237 => "00010000",
        238 => "00010000",
        239 => "00010000",
        240 => "00010000",
        241 => "00010000",
        242 => "00010000",
        243 => "00010000",
        244 => "00010000",
        245 => "00010000",
        246 => "00010000",
        247 => "00010000",
        248 => "00010000",
        249 => "00010000",
        250 => "00010000",
        251 => "00110100",
        252 => "11011111",
        253 => "11011011",
        254 => "00000001",
        255 => "00000001",
        256 => "11011111",
        257 => "10111110",
        258 => "00001100",
        259 => "00010000",
        260 => "00010000",
        261 => "00010100",
        262 => "00010000",
        263 => "00010000",
        264 => "00010000",
        265 => "00010000",
        266 => "00010000",
        267 => "00010000",
        268 => "00010000",
        269 => "00010000",
        270 => "00010000",
        271 => "00010000",
        272 => "00010000",
        273 => "00010000",
        274 => "00010000",
        275 => "00010000",
        276 => "00010000",
        277 => "00010000",
        278 => "00010000",
        279 => "00010000",
        280 => "00010000",
        281 => "00010000",
        282 => "00010000",
        283 => "00010000",
        284 => "00010000",
        285 => "00010000",
        286 => "00010000",
        287 => "00010000",
        288 => "00010000",
        289 => "00010000",
        290 => "00010000",
        291 => "00010000",
        292 => "00010000",
        293 => "00010000",
        294 => "00010000",
        295 => "00010000",
        296 => "00010000",
        297 => "00010000",
        298 => "00010000",
        299 => "00010000",
        300 => "00010000",
        301 => "00010000",
        302 => "00010000",
        303 => "11011111",
        304 => "11011011",
        305 => "00000000",
        306 => "00000001",
        307 => "11011111",
        308 => "10111110",
        309 => "00010000",
        310 => "00010000",
        311 => "00010000",
        312 => "00010000",
        313 => "00010000",
        314 => "00010000",
        315 => "00010000",
        316 => "00010000",
        317 => "00010000",
        318 => "00010000",
        319 => "00010000",
        320 => "00010000",
        321 => "00010000",
        322 => "00010000",
        323 => "00010000",
        324 => "00010000",
        325 => "00010000",
        326 => "00010000",
        327 => "00010000",
        328 => "00010000",
        329 => "00010000",
        330 => "00010000",
        331 => "00010000",
        332 => "00010000",
        333 => "00010000",
        334 => "00010000",
        335 => "00010000",
        336 => "00010000",
        337 => "00010000",
        338 => "00010000",
        339 => "00010000",
        340 => "00010000",
        341 => "00010000",
        342 => "00010000",
        343 => "00010000",
        344 => "00010000",
        345 => "00010000",
        346 => "00010000",
        347 => "00010000",
        348 => "00010000",
        349 => "00010000",
        350 => "00010000",
        351 => "00010000",
        352 => "00010000",
        353 => "00110000",
        354 => "11011111",
        355 => "11011011",
        356 => "00000001",
        357 => "00000001",
        358 => "11011111",
        359 => "10111110",
        360 => "00010000",
        361 => "00010000",
        362 => "00010100",
        363 => "00010000",
        364 => "00010100",
        365 => "00010000",
        366 => "00010000",
        367 => "00010000",
        368 => "00010000",
        369 => "00010000",
        370 => "00010000",
        371 => "00010000",
        372 => "00010000",
        373 => "00010000",
        374 => "00010000",
        375 => "00010000",
        376 => "00010000",
        377 => "00010000",
        378 => "00010000",
        379 => "00010000",
        380 => "00010000",
        381 => "00010000",
        382 => "00010000",
        383 => "00010000",
        384 => "00010000",
        385 => "00010000",
        386 => "00010000",
        387 => "00010000",
        388 => "00010000",
        389 => "00010000",
        390 => "00010000",
        391 => "00010000",
        392 => "00010000",
        393 => "00010000",
        394 => "00010000",
        395 => "00010000",
        396 => "00010000",
        397 => "00010000",
        398 => "00010000",
        399 => "00010000",
        400 => "00010000",
        401 => "00010000",
        402 => "00010000",
        403 => "00010000",
        404 => "00010000",
        405 => "11011111",
        406 => "11011011",
        407 => "00000000",
        408 => "00000000",
        409 => "11011111",
        410 => "10111110",
        411 => "00010000",
        412 => "00010000",
        413 => "00010000",
        414 => "00010000",
        415 => "00010000",
        416 => "00010000",
        417 => "00010000",
        418 => "00010000",
        419 => "00010000",
        420 => "00010000",
        421 => "00010100",
        422 => "00010000",
        423 => "00010000",
        424 => "00010000",
        425 => "00010000",
        426 => "00010000",
        427 => "00010000",
        428 => "00010000",
        429 => "00010000",
        430 => "00010000",
        431 => "00010000",
        432 => "00010000",
        433 => "00010000",
        434 => "00010000",
        435 => "00010000",
        436 => "00010000",
        437 => "00010000",
        438 => "00010000",
        439 => "00010000",
        440 => "00010000",
        441 => "00010000",
        442 => "00010000",
        443 => "00010000",
        444 => "00010000",
        445 => "00010000",
        446 => "00010000",
        447 => "00010000",
        448 => "00010000",
        449 => "00010000",
        450 => "00010000",
        451 => "00010000",
        452 => "00010000",
        453 => "00010000",
        454 => "00010000",
        455 => "00110000",
        456 => "11011111",
        457 => "11011011",
        458 => "00000001",
        459 => "00000000",
        460 => "11111111",
        461 => "10111110",
        462 => "00010000",
        463 => "00010000",
        464 => "00010000",
        465 => "00010000",
        466 => "00010000",
        467 => "00010000",
        468 => "00010000",
        469 => "00010000",
        470 => "00010100",
        471 => "00010000",
        472 => "00010000",
        473 => "00010000",
        474 => "00010000",
        475 => "00010000",
        476 => "00010000",
        477 => "00010000",
        478 => "00010000",
        479 => "00010000",
        480 => "00010000",
        481 => "00010000",
        482 => "00010000",
        483 => "00010000",
        484 => "00010000",
        485 => "00010000",
        486 => "00010100",
        487 => "00010000",
        488 => "00010000",
        489 => "00010000",
        490 => "00010000",
        491 => "00010000",
        492 => "00010000",
        493 => "00010000",
        494 => "00010000",
        495 => "00010000",
        496 => "00010100",
        497 => "00010000",
        498 => "00010000",
        499 => "00010000",
        500 => "00010000",
        501 => "00010000",
        502 => "00010000",
        503 => "00010000",
        504 => "00010000",
        505 => "00010000",
        506 => "00010000",
        507 => "11011111",
        508 => "11011011",
        509 => "00000001",
        510 => "00000001",
        511 => "11111111",
        512 => "10111110",
        513 => "00010000",
        514 => "00010000",
        515 => "00010000",
        516 => "00010000",
        517 => "00010000",
        518 => "00010000",
        519 => "00010000",
        520 => "00010000",
        521 => "00010000",
        522 => "00010000",
        523 => "00010000",
        524 => "00010000",
        525 => "00010000",
        526 => "00010000",
        527 => "00010000",
        528 => "00010000",
        529 => "00010100",
        530 => "00010000",
        531 => "00010000",
        532 => "00010000",
        533 => "00010000",
        534 => "00010000",
        535 => "00010000",
        536 => "00010000",
        537 => "00010100",
        538 => "00010000",
        539 => "00010000",
        540 => "00010000",
        541 => "00010000",
        542 => "00010000",
        543 => "00010000",
        544 => "00010000",
        545 => "00010000",
        546 => "00010000",
        547 => "00010000",
        548 => "00010000",
        549 => "00010100",
        550 => "00010000",
        551 => "00010000",
        552 => "00010000",
        553 => "00010000",
        554 => "00010000",
        555 => "00010000",
        556 => "00010000",
        557 => "00010000",
        558 => "11011111",
        559 => "11011011",
        560 => "00000001",
        561 => "00000001",
        562 => "11111111",
        563 => "10111110",
        564 => "00010000",
        565 => "00010000",
        566 => "00010000",
        567 => "00010000",
        568 => "00010000",
        569 => "00010000",
        570 => "00010100",
        571 => "00010000",
        572 => "00010000",
        573 => "00010000",
        574 => "00010000",
        575 => "00010000",
        576 => "00010000",
        577 => "00010000",
        578 => "00010000",
        579 => "00010000",
        580 => "00010000",
        581 => "00010000",
        582 => "00010000",
        583 => "00110000",
        584 => "00010000",
        585 => "00010000",
        586 => "00010000",
        587 => "00010000",
        588 => "00010000",
        589 => "00010000",
        590 => "00010000",
        591 => "00010000",
        592 => "00010000",
        593 => "00010000",
        594 => "00010000",
        595 => "00010000",
        596 => "00010000",
        597 => "00010000",
        598 => "00010000",
        599 => "00010000",
        600 => "00010000",
        601 => "00010000",
        602 => "00010000",
        603 => "00010000",
        604 => "00010000",
        605 => "00010000",
        606 => "00010000",
        607 => "00010000",
        608 => "00010000",
        609 => "11011111",
        610 => "11011011",
        611 => "00000001",
        612 => "00000001",
        613 => "11011111",
        614 => "10111110",
        615 => "00010000",
        616 => "00010000",
        617 => "00010000",
        618 => "00010000",
        619 => "00010000",
        620 => "00010000",
        621 => "00010000",
        622 => "00010000",
        623 => "00010000",
        624 => "00010000",
        625 => "00010000",
        626 => "00010000",
        627 => "00010000",
        628 => "00010000",
        629 => "00010000",
        630 => "00010000",
        631 => "00010000",
        632 => "00010100",
        633 => "10011101",
        634 => "10111101",
        635 => "01010100",
        636 => "00010000",
        637 => "00010000",
        638 => "00010000",
        639 => "00010000",
        640 => "00010000",
        641 => "00010000",
        642 => "00010000",
        643 => "00010000",
        644 => "00010000",
        645 => "00010000",
        646 => "00010000",
        647 => "00010000",
        648 => "00010000",
        649 => "00010000",
        650 => "00010000",
        651 => "00010000",
        652 => "00010000",
        653 => "00010000",
        654 => "00010100",
        655 => "00010000",
        656 => "00010000",
        657 => "00010000",
        658 => "00010000",
        659 => "00010000",
        660 => "11011111",
        661 => "11011011",
        662 => "00000001",
        663 => "00000001",
        664 => "11011111",
        665 => "10111110",
        666 => "00010000",
        667 => "00010000",
        668 => "00010000",
        669 => "00010000",
        670 => "00010000",
        671 => "00010000",
        672 => "00010000",
        673 => "00010100",
        674 => "00111001",
        675 => "10111110",
        676 => "01111001",
        677 => "00010000",
        678 => "00010000",
        679 => "01010101",
        680 => "10111110",
        681 => "01111101",
        682 => "00001100",
        683 => "00010000",
        684 => "10011110",
        685 => "10111101",
        686 => "01010000",
        687 => "00010000",
        688 => "00010000",
        689 => "00010000",
        690 => "00010000",
        691 => "00010000",
        692 => "00010000",
        693 => "00010000",
        694 => "00010000",
        695 => "00010000",
        696 => "00010000",
        697 => "00010000",
        698 => "00010000",
        699 => "00010000",
        700 => "00010000",
        701 => "00010000",
        702 => "00010000",
        703 => "00010000",
        704 => "00010000",
        705 => "00010000",
        706 => "00010000",
        707 => "00010000",
        708 => "00010000",
        709 => "00010000",
        710 => "00010000",
        711 => "11011111",
        712 => "11011011",
        713 => "00000001",
        714 => "00000001",
        715 => "11011111",
        716 => "10111110",
        717 => "00010000",
        718 => "00010000",
        719 => "00010000",
        720 => "00010000",
        721 => "00010000",
        722 => "00010000",
        723 => "00010000",
        724 => "00010000",
        725 => "00010100",
        726 => "10111110",
        727 => "10111110",
        728 => "00010000",
        729 => "00110000",
        730 => "10011110",
        731 => "10111110",
        732 => "01011000",
        733 => "00010000",
        734 => "00110000",
        735 => "00101100",
        736 => "00110000",
        737 => "00010000",
        738 => "00010000",
        739 => "00010000",
        740 => "00010000",
        741 => "00010000",
        742 => "00010000",
        743 => "00010000",
        744 => "00110000",
        745 => "00010000",
        746 => "00010000",
        747 => "00010000",
        748 => "00010000",
        749 => "00010000",
        750 => "00010000",
        751 => "00010000",
        752 => "00010000",
        753 => "00010000",
        754 => "00010000",
        755 => "00010000",
        756 => "00010000",
        757 => "00010000",
        758 => "00010000",
        759 => "00010000",
        760 => "00010000",
        761 => "00110000",
        762 => "11011111",
        763 => "11011011",
        764 => "00000001",
        765 => "00000001",
        766 => "11011111",
        767 => "10111110",
        768 => "00010000",
        769 => "00010000",
        770 => "00010000",
        771 => "00010000",
        772 => "00010000",
        773 => "00010000",
        774 => "00010000",
        775 => "00010000",
        776 => "00010000",
        777 => "10011110",
        778 => "10111110",
        779 => "01010101",
        780 => "00110000",
        781 => "10111110",
        782 => "10111110",
        783 => "00110100",
        784 => "01011000",
        785 => "10111110",
        786 => "10111110",
        787 => "10111110",
        788 => "01010100",
        789 => "00010000",
        790 => "00010000",
        791 => "00010000",
        792 => "01011001",
        793 => "10111110",
        794 => "10111110",
        795 => "10111110",
        796 => "10011110",
        797 => "01010100",
        798 => "10011110",
        799 => "01011000",
        800 => "00010000",
        801 => "00010000",
        802 => "00010000",
        803 => "01111101",
        804 => "10011101",
        805 => "00010100",
        806 => "00010000",
        807 => "00010000",
        808 => "00010000",
        809 => "00010000",
        810 => "00010000",
        811 => "00010000",
        812 => "00110000",
        813 => "11011111",
        814 => "11011011",
        815 => "00000001",
        816 => "00000001",
        817 => "11011111",
        818 => "10111110",
        819 => "00010000",
        820 => "00010000",
        821 => "00010000",
        822 => "00010000",
        823 => "00010000",
        824 => "00010000",
        825 => "00010000",
        826 => "00010000",
        827 => "00010000",
        828 => "01111110",
        829 => "10111111",
        830 => "01111010",
        831 => "01010001",
        832 => "11011110",
        833 => "10011001",
        834 => "00010000",
        835 => "00010000",
        836 => "00010000",
        837 => "10011101",
        838 => "11011110",
        839 => "01010000",
        840 => "00010000",
        841 => "00010000",
        842 => "00111001",
        843 => "10111110",
        844 => "10011001",
        845 => "01001100",
        846 => "01110101",
        847 => "10111111",
        848 => "10011110",
        849 => "10111110",
        850 => "10011101",
        851 => "00110000",
        852 => "00110000",
        853 => "00110000",
        854 => "10011101",
        855 => "10011101",
        856 => "00010000",
        857 => "00010000",
        858 => "00010000",
        859 => "00010000",
        860 => "00010000",
        861 => "00010000",
        862 => "00010000",
        863 => "00010000",
        864 => "11011111",
        865 => "11011011",
        866 => "00000001",
        867 => "00000000",
        868 => "11011111",
        869 => "10111110",
        870 => "00010000",
        871 => "00010000",
        872 => "00010000",
        873 => "00010000",
        874 => "00010000",
        875 => "00010000",
        876 => "00010000",
        877 => "00010000",
        878 => "00010000",
        879 => "00110101",
        880 => "10111111",
        881 => "10011010",
        882 => "01110101",
        883 => "11011110",
        884 => "01110100",
        885 => "00010000",
        886 => "00010000",
        887 => "00010000",
        888 => "01111101",
        889 => "11011110",
        890 => "01110000",
        891 => "00010000",
        892 => "00010000",
        893 => "01111110",
        894 => "10111111",
        895 => "11011110",
        896 => "11011110",
        897 => "10111110",
        898 => "10111110",
        899 => "10011010",
        900 => "10111110",
        901 => "10011110",
        902 => "01110101",
        903 => "11011110",
        904 => "10011001",
        905 => "11011110",
        906 => "10011001",
        907 => "00010000",
        908 => "00010000",
        909 => "00010000",
        910 => "00010000",
        911 => "00010000",
        912 => "00010000",
        913 => "00010000",
        914 => "00010000",
        915 => "11011111",
        916 => "11011011",
        917 => "00000001",
        918 => "00000000",
        919 => "11011111",
        920 => "10111110",
        921 => "00010000",
        922 => "00010000",
        923 => "00010000",
        924 => "00010000",
        925 => "00010000",
        926 => "00010000",
        927 => "00010000",
        928 => "00010000",
        929 => "00010000",
        930 => "00010000",
        931 => "10111111",
        932 => "11011111",
        933 => "11011110",
        934 => "10111101",
        935 => "00110000",
        936 => "00010000",
        937 => "00010000",
        938 => "00010000",
        939 => "01111110",
        940 => "11011110",
        941 => "01110000",
        942 => "00010000",
        943 => "00010000",
        944 => "10011010",
        945 => "10111110",
        946 => "01111001",
        947 => "00110000",
        948 => "00010000",
        949 => "00001100",
        950 => "00010000",
        951 => "10011110",
        952 => "10111110",
        953 => "10111010",
        954 => "11011110",
        955 => "11011110",
        956 => "11011110",
        957 => "01111001",
        958 => "00010000",
        959 => "00010000",
        960 => "00010000",
        961 => "00010000",
        962 => "00010000",
        963 => "00010000",
        964 => "00010000",
        965 => "00110000",
        966 => "11011111",
        967 => "11011011",
        968 => "00000001",
        969 => "00000000",
        970 => "11011111",
        971 => "10111110",
        972 => "00010000",
        973 => "00010000",
        974 => "00010000",
        975 => "00010000",
        976 => "00010000",
        977 => "00010000",
        978 => "00010000",
        979 => "00010000",
        980 => "00010000",
        981 => "00010000",
        982 => "01111010",
        983 => "11011111",
        984 => "11011110",
        985 => "10011101",
        986 => "00010000",
        987 => "00010000",
        988 => "00010000",
        989 => "00010100",
        990 => "10011110",
        991 => "10111110",
        992 => "01110100",
        993 => "00110000",
        994 => "00010000",
        995 => "01010101",
        996 => "10111110",
        997 => "10011101",
        998 => "00010000",
        999 => "00010000",
        1000 => "00010000",
        1001 => "00010000",
        1002 => "01111110",
        1003 => "10111110",
        1004 => "11011110",
        1005 => "10010101",
        1006 => "11011110",
        1007 => "11011110",
        1008 => "01110100",
        1009 => "00010000",
        1010 => "00010000",
        1011 => "00010000",
        1012 => "00010000",
        1013 => "00010000",
        1014 => "00010000",
        1015 => "00010000",
        1016 => "00110000",
        1017 => "11011111",
        1018 => "11011011",
        1019 => "00000001",
        1020 => "00000001",
        1021 => "11011111",
        1022 => "10111110",
        1023 => "00010000",
        1024 => "00010000",
        1025 => "00010000",
        1026 => "00010000",
        1027 => "00010000",
        1028 => "00010000",
        1029 => "00010000",
        1030 => "00010000",
        1031 => "00010000",
        1032 => "00010000",
        1033 => "01010101",
        1034 => "10111110",
        1035 => "10111110",
        1036 => "01011000",
        1037 => "00010000",
        1038 => "00010100",
        1039 => "01111101",
        1040 => "10111110",
        1041 => "10111110",
        1042 => "10111110",
        1043 => "10111110",
        1044 => "10011101",
        1045 => "00110100",
        1046 => "00010000",
        1047 => "01011001",
        1048 => "10111110",
        1049 => "10111110",
        1050 => "10011110",
        1051 => "10011101",
        1052 => "00110100",
        1053 => "01011001",
        1054 => "10111110",
        1055 => "10011101",
        1056 => "00110000",
        1057 => "10011101",
        1058 => "10111101",
        1059 => "00110100",
        1060 => "00010000",
        1061 => "00010000",
        1062 => "00010000",
        1063 => "00010000",
        1064 => "00010000",
        1065 => "00010000",
        1066 => "00010000",
        1067 => "00110000",
        1068 => "11011111",
        1069 => "11011011",
        1070 => "00000001",
        1071 => "00000001",
        1072 => "11011111",
        1073 => "10111110",
        1074 => "00010000",
        1075 => "00010000",
        1076 => "00010000",
        1077 => "00010000",
        1078 => "00010000",
        1079 => "00010000",
        1080 => "00010000",
        1081 => "00010000",
        1082 => "00010100",
        1083 => "00010000",
        1084 => "00010000",
        1085 => "00010000",
        1086 => "00010000",
        1087 => "00010000",
        1088 => "00010000",
        1089 => "00010000",
        1090 => "00010000",
        1091 => "00010000",
        1092 => "00010000",
        1093 => "00001100",
        1094 => "00010000",
        1095 => "00010000",
        1096 => "00010000",
        1097 => "00010000",
        1098 => "00010000",
        1099 => "00010000",
        1100 => "00010000",
        1101 => "00010000",
        1102 => "00010000",
        1103 => "00010000",
        1104 => "00010000",
        1105 => "00010000",
        1106 => "00001100",
        1107 => "00010000",
        1108 => "00010000",
        1109 => "00010000",
        1110 => "00010000",
        1111 => "00010000",
        1112 => "00010000",
        1113 => "00010000",
        1114 => "00010000",
        1115 => "00010000",
        1116 => "00010000",
        1117 => "00010000",
        1118 => "00110000",
        1119 => "11011111",
        1120 => "11011011",
        1121 => "00000001",
        1122 => "00000001",
        1123 => "11011111",
        1124 => "10111110",
        1125 => "00010000",
        1126 => "00010000",
        1127 => "00010000",
        1128 => "00010100",
        1129 => "00010000",
        1130 => "00010000",
        1131 => "00010000",
        1132 => "00010000",
        1133 => "00010100",
        1134 => "00010000",
        1135 => "00010000",
        1136 => "00010000",
        1137 => "00010000",
        1138 => "00010000",
        1139 => "00010000",
        1140 => "00010000",
        1141 => "00010000",
        1142 => "00010000",
        1143 => "00010000",
        1144 => "00010000",
        1145 => "00010000",
        1146 => "00010000",
        1147 => "00010000",
        1148 => "00010000",
        1149 => "00010000",
        1150 => "00010000",
        1151 => "00010000",
        1152 => "00010000",
        1153 => "00010000",
        1154 => "00010000",
        1155 => "00010000",
        1156 => "00010000",
        1157 => "00010100",
        1158 => "00010000",
        1159 => "00010000",
        1160 => "00010000",
        1161 => "00010000",
        1162 => "00010000",
        1163 => "00010000",
        1164 => "00010000",
        1165 => "00010000",
        1166 => "00010000",
        1167 => "00010000",
        1168 => "00010000",
        1169 => "00110000",
        1170 => "11011111",
        1171 => "11011011",
        1172 => "00000001",
        1173 => "00000001",
        1174 => "11011111",
        1175 => "10111110",
        1176 => "00010000",
        1177 => "00010000",
        1178 => "00010000",
        1179 => "00010000",
        1180 => "00010000",
        1181 => "00010000",
        1182 => "00010000",
        1183 => "00010000",
        1184 => "00010000",
        1185 => "00010000",
        1186 => "00010000",
        1187 => "00010000",
        1188 => "00010000",
        1189 => "00010000",
        1190 => "00010000",
        1191 => "00010000",
        1192 => "00010000",
        1193 => "00010000",
        1194 => "00010100",
        1195 => "00010000",
        1196 => "00010000",
        1197 => "00010000",
        1198 => "00010000",
        1199 => "00010000",
        1200 => "00010000",
        1201 => "00010000",
        1202 => "00010000",
        1203 => "00010000",
        1204 => "00010000",
        1205 => "00010000",
        1206 => "00010000",
        1207 => "00010000",
        1208 => "00010000",
        1209 => "00010000",
        1210 => "00010000",
        1211 => "00010000",
        1212 => "00010000",
        1213 => "00010000",
        1214 => "00010000",
        1215 => "00010000",
        1216 => "00010000",
        1217 => "00010100",
        1218 => "00010100",
        1219 => "00010000",
        1220 => "00110000",
        1221 => "11011111",
        1222 => "11011011",
        1223 => "00000001",
        1224 => "00000000",
        1225 => "11011111",
        1226 => "10111110",
        1227 => "00010000",
        1228 => "00010000",
        1229 => "00010000",
        1230 => "00010000",
        1231 => "00010000",
        1232 => "00010000",
        1233 => "00010000",
        1234 => "00010000",
        1235 => "00010000",
        1236 => "00010000",
        1237 => "00010000",
        1238 => "00010000",
        1239 => "00010000",
        1240 => "00010000",
        1241 => "00010000",
        1242 => "00010000",
        1243 => "00010000",
        1244 => "00010000",
        1245 => "00010000",
        1246 => "00010000",
        1247 => "00010000",
        1248 => "00010000",
        1249 => "00010000",
        1250 => "00010000",
        1251 => "00010000",
        1252 => "00010000",
        1253 => "00010000",
        1254 => "00010000",
        1255 => "00010000",
        1256 => "00010000",
        1257 => "00010000",
        1258 => "00010000",
        1259 => "00010000",
        1260 => "00010000",
        1261 => "00010000",
        1262 => "00010000",
        1263 => "00010000",
        1264 => "00010100",
        1265 => "00010000",
        1266 => "00010000",
        1267 => "00010000",
        1268 => "00010100",
        1269 => "00010000",
        1270 => "00010000",
        1271 => "00110000",
        1272 => "11011111",
        1273 => "11011011",
        1274 => "00000001",
        1275 => "00000000",
        1276 => "11011111",
        1277 => "10111110",
        1278 => "00010000",
        1279 => "00010000",
        1280 => "00010000",
        1281 => "00010000",
        1282 => "00010000",
        1283 => "00010000",
        1284 => "00010000",
        1285 => "00010000",
        1286 => "00010000",
        1287 => "00010000",
        1288 => "00010000",
        1289 => "00010000",
        1290 => "00010000",
        1291 => "00010000",
        1292 => "00010000",
        1293 => "00010000",
        1294 => "00010000",
        1295 => "00010000",
        1296 => "00010000",
        1297 => "00010000",
        1298 => "00010000",
        1299 => "00010000",
        1300 => "00010000",
        1301 => "00010000",
        1302 => "00010000",
        1303 => "00010000",
        1304 => "00010000",
        1305 => "00010000",
        1306 => "00010000",
        1307 => "00010000",
        1308 => "00010000",
        1309 => "00010000",
        1310 => "00010000",
        1311 => "00010000",
        1312 => "00010000",
        1313 => "00010000",
        1314 => "00010000",
        1315 => "00010000",
        1316 => "00010100",
        1317 => "00010100",
        1318 => "00010000",
        1319 => "00010000",
        1320 => "00010000",
        1321 => "00010000",
        1322 => "00110000",
        1323 => "11011111",
        1324 => "11011011",
        1325 => "00000001",
        1326 => "00100001",
        1327 => "11111111",
        1328 => "10111110",
        1329 => "00010000",
        1330 => "00010000",
        1331 => "00010000",
        1332 => "00010000",
        1333 => "00010000",
        1334 => "00010000",
        1335 => "00010000",
        1336 => "00010000",
        1337 => "00010000",
        1338 => "00010000",
        1339 => "00010000",
        1340 => "00010000",
        1341 => "00010000",
        1342 => "00010000",
        1343 => "00010000",
        1344 => "00010000",
        1345 => "00010000",
        1346 => "00010000",
        1347 => "00010000",
        1348 => "00010000",
        1349 => "00010000",
        1350 => "00010000",
        1351 => "00010000",
        1352 => "00010000",
        1353 => "00010000",
        1354 => "00010000",
        1355 => "00010000",
        1356 => "00010000",
        1357 => "00010000",
        1358 => "00010000",
        1359 => "00010000",
        1360 => "00010000",
        1361 => "00010000",
        1362 => "00010000",
        1363 => "00010000",
        1364 => "00010000",
        1365 => "00010000",
        1366 => "00010000",
        1367 => "00010000",
        1368 => "00010000",
        1369 => "00010000",
        1370 => "00010000",
        1371 => "00010000",
        1372 => "00010000",
        1373 => "00010000",
        1374 => "11011111",
        1375 => "11011011",
        1376 => "00000001",
        1377 => "00100000",
        1378 => "11111111",
        1379 => "10111110",
        1380 => "00010000",
        1381 => "00010000",
        1382 => "00010000",
        1383 => "00010000",
        1384 => "00010000",
        1385 => "00010000",
        1386 => "00010000",
        1387 => "00010000",
        1388 => "00010000",
        1389 => "00010000",
        1390 => "00010000",
        1391 => "00010000",
        1392 => "00010000",
        1393 => "00010000",
        1394 => "00010000",
        1395 => "00010000",
        1396 => "00010000",
        1397 => "00010000",
        1398 => "00010000",
        1399 => "00010000",
        1400 => "00010000",
        1401 => "00010000",
        1402 => "00010000",
        1403 => "00010000",
        1404 => "00010000",
        1405 => "00010000",
        1406 => "00010000",
        1407 => "00010000",
        1408 => "00010000",
        1409 => "00010000",
        1410 => "00010000",
        1411 => "00010000",
        1412 => "00010000",
        1413 => "00010000",
        1414 => "00010000",
        1415 => "00010000",
        1416 => "00010000",
        1417 => "00010000",
        1418 => "00010000",
        1419 => "00010000",
        1420 => "00010000",
        1421 => "00010000",
        1422 => "00010000",
        1423 => "00010000",
        1424 => "00010000",
        1425 => "11011111",
        1426 => "11011011",
        1427 => "00000001",
        1428 => "00000001",
        1429 => "11011111",
        1430 => "10111110",
        1431 => "00001100",
        1432 => "00010000",
        1433 => "00010000",
        1434 => "00010000",
        1435 => "00010000",
        1436 => "00010000",
        1437 => "00010000",
        1438 => "00010000",
        1439 => "00010000",
        1440 => "00010000",
        1441 => "00010000",
        1442 => "00010000",
        1443 => "00010000",
        1444 => "00010000",
        1445 => "00010000",
        1446 => "00010000",
        1447 => "00010000",
        1448 => "00010000",
        1449 => "00010000",
        1450 => "00010000",
        1451 => "00010000",
        1452 => "00010000",
        1453 => "00010000",
        1454 => "00010000",
        1455 => "00010000",
        1456 => "00010000",
        1457 => "00010000",
        1458 => "00010000",
        1459 => "00010000",
        1460 => "00010100",
        1461 => "00010100",
        1462 => "00010000",
        1463 => "00010000",
        1464 => "00010000",
        1465 => "00010000",
        1466 => "00010000",
        1467 => "00010000",
        1468 => "00010000",
        1469 => "00010000",
        1470 => "00010000",
        1471 => "00010000",
        1472 => "00010000",
        1473 => "00010000",
        1474 => "00010000",
        1475 => "00010000",
        1476 => "11011111",
        1477 => "11011011",
        1478 => "00000001",
        1479 => "00000001",
        1480 => "11011111",
        1481 => "10111110",
        1482 => "00110000",
        1483 => "00010000",
        1484 => "00010000",
        1485 => "00010000",
        1486 => "00010000",
        1487 => "00010000",
        1488 => "00010000",
        1489 => "00010000",
        1490 => "00010000",
        1491 => "00010000",
        1492 => "00010000",
        1493 => "00010000",
        1494 => "00010000",
        1495 => "00010000",
        1496 => "00010000",
        1497 => "00010000",
        1498 => "00010000",
        1499 => "00010000",
        1500 => "00010000",
        1501 => "00010000",
        1502 => "00010000",
        1503 => "00010000",
        1504 => "00010000",
        1505 => "00010000",
        1506 => "00010000",
        1507 => "00010000",
        1508 => "00010000",
        1509 => "00010000",
        1510 => "00010000",
        1511 => "00010000",
        1512 => "00010000",
        1513 => "00010000",
        1514 => "00010000",
        1515 => "00010000",
        1516 => "00010000",
        1517 => "00010000",
        1518 => "00010000",
        1519 => "00010000",
        1520 => "00010000",
        1521 => "00010000",
        1522 => "00010000",
        1523 => "00010000",
        1524 => "00010000",
        1525 => "00010000",
        1526 => "01010100",
        1527 => "11011111",
        1528 => "11011011",
        1529 => "00000001",
        1530 => "00000001",
        1531 => "10010111",
        1532 => "11011111",
        1533 => "10010101",
        1534 => "01010000",
        1535 => "00110000",
        1536 => "00010000",
        1537 => "00110000",
        1538 => "00110000",
        1539 => "00110000",
        1540 => "00110000",
        1541 => "00110000",
        1542 => "00110000",
        1543 => "00110000",
        1544 => "00110000",
        1545 => "00110000",
        1546 => "00110000",
        1547 => "00110000",
        1548 => "00110000",
        1549 => "00110000",
        1550 => "00110000",
        1551 => "00110000",
        1552 => "00110000",
        1553 => "00110000",
        1554 => "00110000",
        1555 => "00110000",
        1556 => "00110000",
        1557 => "00010000",
        1558 => "00010000",
        1559 => "00110000",
        1560 => "00110000",
        1561 => "00110000",
        1562 => "00110000",
        1563 => "00110000",
        1564 => "00110000",
        1565 => "00110000",
        1566 => "00110000",
        1567 => "00110000",
        1568 => "00110000",
        1569 => "00110000",
        1570 => "00110000",
        1571 => "00110000",
        1572 => "00110000",
        1573 => "00110000",
        1574 => "00110000",
        1575 => "00110000",
        1576 => "01010100",
        1577 => "10011010",
        1578 => "11011111",
        1579 => "10010010",
        1580 => "00000001",
        1581 => "00000001",
        1582 => "00100101",
        1583 => "11011011",
        1584 => "11011111",
        1585 => "11011111",
        1586 => "11011111",
        1587 => "11011111",
        1588 => "11011111",
        1589 => "11011111",
        1590 => "11011111",
        1591 => "11011111",
        1592 => "11011111",
        1593 => "11011111",
        1594 => "11011111",
        1595 => "11011111",
        1596 => "11011111",
        1597 => "11011111",
        1598 => "11011111",
        1599 => "11011111",
        1600 => "11011111",
        1601 => "11011111",
        1602 => "11011111",
        1603 => "11011111",
        1604 => "11011111",
        1605 => "11011111",
        1606 => "11011111",
        1607 => "11011111",
        1608 => "11011111",
        1609 => "11011111",
        1610 => "11011111",
        1611 => "11011111",
        1612 => "11011111",
        1613 => "11011111",
        1614 => "11011111",
        1615 => "11011111",
        1616 => "11011111",
        1617 => "11011111",
        1618 => "11011111",
        1619 => "11011111",
        1620 => "11011111",
        1621 => "11011111",
        1622 => "11011111",
        1623 => "11011111",
        1624 => "11011111",
        1625 => "11011111",
        1626 => "11011111",
        1627 => "11011111",
        1628 => "11011111",
        1629 => "10111011",
        1630 => "00000001",
        1631 => "00000001",
        1632 => "00000001",
        1633 => "00000001",
        1634 => "00100101",
        1635 => "10010011",
        1636 => "11011011",
        1637 => "11011111",
        1638 => "11011011",
        1639 => "11011111",
        1640 => "11011011",
        1641 => "11011011",
        1642 => "11011011",
        1643 => "11011011",
        1644 => "11011011",
        1645 => "11011011",
        1646 => "11011011",
        1647 => "11011011",
        1648 => "11011011",
        1649 => "11011011",
        1650 => "11011011",
        1651 => "11011011",
        1652 => "11011011",
        1653 => "11011011",
        1654 => "11011011",
        1655 => "11011011",
        1656 => "11011011",
        1657 => "11011011",
        1658 => "11011011",
        1659 => "11011111",
        1660 => "11011011",
        1661 => "11011011",
        1662 => "11011011",
        1663 => "11011011",
        1664 => "11011011",
        1665 => "11011011",
        1666 => "11011011",
        1667 => "11011011",
        1668 => "11011011",
        1669 => "11011011",
        1670 => "11011011",
        1671 => "11011011",
        1672 => "11011111",
        1673 => "11011011",
        1674 => "11011011",
        1675 => "11011011",
        1676 => "11011011",
        1677 => "11011111",
        1678 => "10111011",
        1679 => "10010010",
        1680 => "00000001",
        1681 => "00000001",
        1682 => "00000001",
        1683 => "00000001",
        1684 => "00000001",
        1685 => "00000001",
        1686 => "00000001",
        1687 => "00000000",
        1688 => "00000000",
        1689 => "00000000",
        1690 => "00000000",
        1691 => "00000000",
        1692 => "00000000",
        1693 => "00000000",
        1694 => "00000000",
        1695 => "00000000",
        1696 => "00000000",
        1697 => "00000000",
        1698 => "00000000",
        1699 => "00000000",
        1700 => "00000000",
        1701 => "00000000",
        1702 => "00000000",
        1703 => "00000000",
        1704 => "00000000",
        1705 => "00000000",
        1706 => "00000000",
        1707 => "00000000",
        1708 => "00000000",
        1709 => "00000000",
        1710 => "00000000",
        1711 => "00000000",
        1712 => "00000000",
        1713 => "00000000",
        1714 => "00000000",
        1715 => "00000000",
        1716 => "00000000",
        1717 => "00000000",
        1718 => "00000000",
        1719 => "00000000",
        1720 => "00000000",
        1721 => "00000000",
        1722 => "00000000",
        1723 => "00000000",
        1724 => "00000000",
        1725 => "00000000",
        1726 => "00000000",
        1727 => "00000000",
        1728 => "00000000",
        1729 => "00000000",
        1730 => "00000000",
        1731 => "00000001",
        1732 => "00000001",
        1733 => "00000001");
begin

    process(clk)
    begin
    
        if rising_edge(clk) then
            if rst = '1' then
                view <= (others => (others => '0'));
            else
                dout <= view(to_integer(unsigned(addr)));
            end if;
        end if;
    end process;
end Behavioral;
